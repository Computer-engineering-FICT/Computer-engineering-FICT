* /root/laba15/1.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/1NPN.model

*----------------------------------------------

R_R2 4 2 300 
V_V2 4 0 dc 10 
Q_Q1 2 3 0 1NPN 
R_R1 1 3 2k 
V_V1 1 0 dc 0.0 ac 0.0 PULSE 0.0 5 0 0.01u 0.01u 0.5u 1u 
vtpi@1 1 3 0
*----------------------------------------------

.tran 1e-07 1e-06 0 
.print tran  v(4)
.op

.end
