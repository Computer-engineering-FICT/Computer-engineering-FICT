* /root/laba4/4_2.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/2NMOS.model
*----------------------------------------------

 
M_M1 3 1 2 0 nmos 
V_V2 3 0 dc 10 
V_V1 1 0 dc 0.0 ac 0.0 sin(0.0 5 10000 0 0) 
R_R1 2 0 1000 

*----------------------------------------------

.dc V_V1 0 15 0.01
.print dc   v(1)
.op

.end
