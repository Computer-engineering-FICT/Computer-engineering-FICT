* /root/laba7/2.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/UA741.model

*----------------------------------------------

V_V1 5 0 dc 0 ac 100m sin(0.0 1 10000 0 0) 
R_R3 5 4 1 
V_V2 3 0 dc 10 
R_R2 0 1 10k 
R_R1 1 2 10k 
X_U1 4 1 3 6 2  UA741 
V_V3 0 6 dc 10 
VTPI@1 5 4 0
*----------------------------------------------

.dc V_V1 -10 10 0.1
.print dc   v(0)
.op

.end
