* /root/laba9/4.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/UA741.model

*----------------------------------------------

V_V3 6 0 dc 0.0 ac 100 sin(0.0 10 10000 0 0) 
R_R1 6 1 5k 
V_V1 5 0 dc 5 
R_R2 1 2 10k 
X_U1 3 1 5 7 2 UA741 
V_V2 0 7 dc 5 
C_C2 2 4 1e-8 IC=0 
C_C1 3 0 1e-8 IC=0 
R_R4 4 3 10k 
R_R3 3 0 15k 

*----------------------------------------------

.ac DEC 10 1 1e+08
.print ac  vm(1)
.op

.end
