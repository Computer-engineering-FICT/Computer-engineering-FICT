* /root/laba1/1.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 

*----------------------------------------------

V_V1 1 0 dc 0.0 ac 1.0 sin(0.0 10 10000 0 0) 
R_R1 2 0 100000 
C_C1 1 2 0.59n IC=0 

*----------------------------------------------

.tran 3e-06 0.0003 0 UIC
.print tran  v(2)
.op

.end
