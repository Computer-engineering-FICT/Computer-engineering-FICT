* /root/laba15/3.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/1NPN.model

*----------------------------------------------

R_R4 3 0 1k 
R_R3 3 5 1 
R_R1 2 3 2k 
R_R2 1 4 300 
Q_Q1 4 5 0 1NPN 
V_V1 2 0 dc 0.0 ac 0.0 PULSE 0.0 10 0 0.01u 0.01u 0.5u 1u 
V_V2 1 0 dc 10 
vtpi@1 3 5 0
*----------------------------------------------

.tran 1e-07 5e-06 0 UIC
.print tran  v(1)
.op

.end
