* /root/laba1/3.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 

*----------------------------------------------

R_R1 2 1 1000 
C_C1 1 0 0.59n IC=0 
V_V1 2 0 dc 0.0 ac 0.0 PULSE 0 10 20u 0.5u 0.5u 30u 120u 

*----------------------------------------------

.tran 1e-06 0.0001 0 UIC
.print tran  v(2)
.op

.end
