-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_mux 

-- ============================================================
-- File Name: lpm_mux0.vhd
-- Megafunction Name(s):
-- 			lpm_mux
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 222 10/21/2009 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2009 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY lpm_mux0 IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data0x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data100x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data101x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data102x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data103x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data104x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data105x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data106x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data107x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data108x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data109x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data110x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data111x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data112x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data113x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data114x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data115x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data116x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data117x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data118x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data119x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data120x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data121x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data122x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data123x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data124x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data125x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data126x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data127x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data128x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data129x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data130x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data131x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data132x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data133x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data134x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data135x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data136x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data137x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data138x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data139x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data140x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data141x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data142x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data143x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data144x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data145x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data146x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data147x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data148x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data149x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data150x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data151x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data152x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data153x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data154x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data155x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data156x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data157x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data158x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data159x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data160x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data161x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data162x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data163x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data164x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data165x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data166x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data167x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data168x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data169x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data16x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data170x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data171x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data172x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data173x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data174x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data175x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data176x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data177x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data178x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data179x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data17x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data180x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data181x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data182x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data183x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data184x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data185x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data186x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data187x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data188x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data189x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data18x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data190x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data191x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data192x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data193x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data194x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data195x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data196x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data197x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data198x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data199x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data19x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data200x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data201x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data202x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data203x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data204x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data205x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data206x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data207x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data208x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data209x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data20x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data210x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data211x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data212x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data213x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data214x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data215x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data216x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data217x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data218x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data219x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data21x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data220x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data221x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data222x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data223x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data224x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data225x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data226x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data227x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data228x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data229x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data22x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data230x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data231x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data232x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data233x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data234x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data235x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data236x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data237x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data238x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data239x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data23x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data240x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data241x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data242x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data243x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data244x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data245x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data246x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data247x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data248x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data249x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data24x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data250x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data251x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data252x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data253x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data254x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data255x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data25x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data26x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data27x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data28x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data29x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data30x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data31x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data32x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data33x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data34x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data35x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data36x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data37x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data38x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data39x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data40x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data41x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data42x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data43x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data44x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data45x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data46x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data47x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data48x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data49x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data50x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data51x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data52x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data53x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data54x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data55x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data56x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data57x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data58x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data59x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data60x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data61x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data62x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data63x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data64x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data65x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data66x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data67x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data68x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data69x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data70x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data71x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data72x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data73x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data74x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data75x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data76x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data77x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data78x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data79x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data80x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data81x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data82x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data83x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data84x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data85x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data86x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data87x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data88x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data89x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data90x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data91x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data92x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data93x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data94x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data95x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data96x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data97x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data98x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data99x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (39 DOWNTO 0)
	);
END lpm_mux0;


ARCHITECTURE SYN OF lpm_mux0 IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_2D (255 DOWNTO 0, 39 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire19	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire20	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire21	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire22	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire23	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire24	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire25	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire26	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire27	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire28	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire29	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire30	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire31	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire32	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire33	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire34	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire35	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire36	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire37	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire38	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire39	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire40	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire41	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire42	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire43	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire44	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire45	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire46	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire47	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire48	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire49	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire50	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire51	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire52	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire53	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire54	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire55	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire56	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire57	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire58	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire59	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire60	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire61	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire62	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire63	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire64	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire65	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire66	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire67	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire68	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire69	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire70	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire71	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire72	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire73	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire74	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire75	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire76	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire77	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire78	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire79	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire80	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire81	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire82	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire83	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire84	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire85	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire86	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire87	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire88	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire89	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire90	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire91	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire92	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire93	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire94	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire95	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire96	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire97	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire98	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire99	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire100	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire101	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire102	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire103	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire104	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire105	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire106	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire107	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire108	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire109	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire110	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire111	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire112	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire113	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire114	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire115	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire116	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire117	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire118	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire119	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire120	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire121	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire122	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire123	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire124	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire125	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire126	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire127	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire128	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire129	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire130	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire131	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire132	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire133	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire134	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire135	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire136	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire137	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire138	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire139	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire140	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire141	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire142	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire143	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire144	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire145	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire146	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire147	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire148	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire149	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire150	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire151	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire152	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire153	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire154	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire155	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire156	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire157	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire158	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire159	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire160	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire161	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire162	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire163	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire164	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire165	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire166	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire167	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire168	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire169	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire170	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire171	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire172	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire173	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire174	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire175	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire176	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire177	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire178	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire179	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire180	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire181	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire182	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire183	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire184	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire185	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire186	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire187	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire188	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire189	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire190	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire191	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire192	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire193	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire194	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire195	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire196	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire197	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire198	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire199	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire200	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire201	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire202	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire203	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire204	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire205	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire206	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire207	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire208	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire209	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire210	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire211	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire212	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire213	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire214	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire215	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire216	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire217	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire218	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire219	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire220	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire221	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire222	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire223	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire224	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire225	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire226	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire227	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire228	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire229	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire230	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire231	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire232	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire233	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire234	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire235	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire236	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire237	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire238	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire239	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire240	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire241	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire242	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire243	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire244	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire245	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire246	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire247	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire248	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire249	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire250	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire251	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire252	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire253	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire254	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire255	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire256	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire257	: STD_LOGIC_VECTOR (39 DOWNTO 0);

BEGIN
	sub_wire257    <= data0x(39 DOWNTO 0);
	sub_wire256    <= data1x(39 DOWNTO 0);
	sub_wire255    <= data2x(39 DOWNTO 0);
	sub_wire254    <= data3x(39 DOWNTO 0);
	sub_wire253    <= data4x(39 DOWNTO 0);
	sub_wire252    <= data5x(39 DOWNTO 0);
	sub_wire251    <= data6x(39 DOWNTO 0);
	sub_wire250    <= data7x(39 DOWNTO 0);
	sub_wire249    <= data8x(39 DOWNTO 0);
	sub_wire248    <= data9x(39 DOWNTO 0);
	sub_wire247    <= data10x(39 DOWNTO 0);
	sub_wire246    <= data11x(39 DOWNTO 0);
	sub_wire245    <= data12x(39 DOWNTO 0);
	sub_wire244    <= data13x(39 DOWNTO 0);
	sub_wire243    <= data14x(39 DOWNTO 0);
	sub_wire242    <= data15x(39 DOWNTO 0);
	sub_wire241    <= data16x(39 DOWNTO 0);
	sub_wire240    <= data17x(39 DOWNTO 0);
	sub_wire239    <= data18x(39 DOWNTO 0);
	sub_wire238    <= data19x(39 DOWNTO 0);
	sub_wire237    <= data20x(39 DOWNTO 0);
	sub_wire236    <= data21x(39 DOWNTO 0);
	sub_wire235    <= data22x(39 DOWNTO 0);
	sub_wire234    <= data23x(39 DOWNTO 0);
	sub_wire233    <= data24x(39 DOWNTO 0);
	sub_wire232    <= data25x(39 DOWNTO 0);
	sub_wire231    <= data26x(39 DOWNTO 0);
	sub_wire230    <= data27x(39 DOWNTO 0);
	sub_wire229    <= data28x(39 DOWNTO 0);
	sub_wire228    <= data29x(39 DOWNTO 0);
	sub_wire227    <= data30x(39 DOWNTO 0);
	sub_wire226    <= data31x(39 DOWNTO 0);
	sub_wire225    <= data32x(39 DOWNTO 0);
	sub_wire224    <= data33x(39 DOWNTO 0);
	sub_wire223    <= data34x(39 DOWNTO 0);
	sub_wire222    <= data35x(39 DOWNTO 0);
	sub_wire221    <= data36x(39 DOWNTO 0);
	sub_wire220    <= data37x(39 DOWNTO 0);
	sub_wire219    <= data38x(39 DOWNTO 0);
	sub_wire218    <= data39x(39 DOWNTO 0);
	sub_wire217    <= data40x(39 DOWNTO 0);
	sub_wire216    <= data41x(39 DOWNTO 0);
	sub_wire215    <= data42x(39 DOWNTO 0);
	sub_wire214    <= data43x(39 DOWNTO 0);
	sub_wire213    <= data44x(39 DOWNTO 0);
	sub_wire212    <= data45x(39 DOWNTO 0);
	sub_wire211    <= data46x(39 DOWNTO 0);
	sub_wire210    <= data47x(39 DOWNTO 0);
	sub_wire209    <= data48x(39 DOWNTO 0);
	sub_wire208    <= data49x(39 DOWNTO 0);
	sub_wire207    <= data50x(39 DOWNTO 0);
	sub_wire206    <= data51x(39 DOWNTO 0);
	sub_wire205    <= data52x(39 DOWNTO 0);
	sub_wire204    <= data53x(39 DOWNTO 0);
	sub_wire203    <= data54x(39 DOWNTO 0);
	sub_wire202    <= data55x(39 DOWNTO 0);
	sub_wire201    <= data56x(39 DOWNTO 0);
	sub_wire200    <= data57x(39 DOWNTO 0);
	sub_wire199    <= data58x(39 DOWNTO 0);
	sub_wire198    <= data59x(39 DOWNTO 0);
	sub_wire197    <= data60x(39 DOWNTO 0);
	sub_wire196    <= data61x(39 DOWNTO 0);
	sub_wire195    <= data62x(39 DOWNTO 0);
	sub_wire194    <= data63x(39 DOWNTO 0);
	sub_wire193    <= data64x(39 DOWNTO 0);
	sub_wire192    <= data65x(39 DOWNTO 0);
	sub_wire191    <= data66x(39 DOWNTO 0);
	sub_wire190    <= data67x(39 DOWNTO 0);
	sub_wire189    <= data68x(39 DOWNTO 0);
	sub_wire188    <= data69x(39 DOWNTO 0);
	sub_wire187    <= data70x(39 DOWNTO 0);
	sub_wire186    <= data71x(39 DOWNTO 0);
	sub_wire185    <= data72x(39 DOWNTO 0);
	sub_wire184    <= data73x(39 DOWNTO 0);
	sub_wire183    <= data74x(39 DOWNTO 0);
	sub_wire182    <= data75x(39 DOWNTO 0);
	sub_wire181    <= data76x(39 DOWNTO 0);
	sub_wire180    <= data77x(39 DOWNTO 0);
	sub_wire179    <= data78x(39 DOWNTO 0);
	sub_wire178    <= data79x(39 DOWNTO 0);
	sub_wire177    <= data80x(39 DOWNTO 0);
	sub_wire176    <= data81x(39 DOWNTO 0);
	sub_wire175    <= data82x(39 DOWNTO 0);
	sub_wire174    <= data83x(39 DOWNTO 0);
	sub_wire173    <= data84x(39 DOWNTO 0);
	sub_wire172    <= data85x(39 DOWNTO 0);
	sub_wire171    <= data86x(39 DOWNTO 0);
	sub_wire170    <= data87x(39 DOWNTO 0);
	sub_wire169    <= data88x(39 DOWNTO 0);
	sub_wire168    <= data89x(39 DOWNTO 0);
	sub_wire167    <= data90x(39 DOWNTO 0);
	sub_wire166    <= data91x(39 DOWNTO 0);
	sub_wire165    <= data92x(39 DOWNTO 0);
	sub_wire164    <= data93x(39 DOWNTO 0);
	sub_wire163    <= data94x(39 DOWNTO 0);
	sub_wire162    <= data95x(39 DOWNTO 0);
	sub_wire161    <= data96x(39 DOWNTO 0);
	sub_wire160    <= data97x(39 DOWNTO 0);
	sub_wire159    <= data98x(39 DOWNTO 0);
	sub_wire158    <= data99x(39 DOWNTO 0);
	sub_wire157    <= data100x(39 DOWNTO 0);
	sub_wire156    <= data101x(39 DOWNTO 0);
	sub_wire155    <= data102x(39 DOWNTO 0);
	sub_wire154    <= data103x(39 DOWNTO 0);
	sub_wire153    <= data104x(39 DOWNTO 0);
	sub_wire152    <= data105x(39 DOWNTO 0);
	sub_wire151    <= data106x(39 DOWNTO 0);
	sub_wire150    <= data107x(39 DOWNTO 0);
	sub_wire149    <= data108x(39 DOWNTO 0);
	sub_wire148    <= data109x(39 DOWNTO 0);
	sub_wire147    <= data110x(39 DOWNTO 0);
	sub_wire146    <= data111x(39 DOWNTO 0);
	sub_wire145    <= data112x(39 DOWNTO 0);
	sub_wire144    <= data113x(39 DOWNTO 0);
	sub_wire143    <= data114x(39 DOWNTO 0);
	sub_wire142    <= data115x(39 DOWNTO 0);
	sub_wire141    <= data116x(39 DOWNTO 0);
	sub_wire140    <= data117x(39 DOWNTO 0);
	sub_wire139    <= data118x(39 DOWNTO 0);
	sub_wire138    <= data119x(39 DOWNTO 0);
	sub_wire137    <= data120x(39 DOWNTO 0);
	sub_wire136    <= data121x(39 DOWNTO 0);
	sub_wire135    <= data122x(39 DOWNTO 0);
	sub_wire134    <= data123x(39 DOWNTO 0);
	sub_wire133    <= data124x(39 DOWNTO 0);
	sub_wire132    <= data125x(39 DOWNTO 0);
	sub_wire131    <= data126x(39 DOWNTO 0);
	sub_wire130    <= data127x(39 DOWNTO 0);
	sub_wire129    <= data128x(39 DOWNTO 0);
	sub_wire128    <= data129x(39 DOWNTO 0);
	sub_wire127    <= data130x(39 DOWNTO 0);
	sub_wire126    <= data131x(39 DOWNTO 0);
	sub_wire125    <= data132x(39 DOWNTO 0);
	sub_wire124    <= data133x(39 DOWNTO 0);
	sub_wire123    <= data134x(39 DOWNTO 0);
	sub_wire122    <= data135x(39 DOWNTO 0);
	sub_wire121    <= data136x(39 DOWNTO 0);
	sub_wire120    <= data137x(39 DOWNTO 0);
	sub_wire119    <= data138x(39 DOWNTO 0);
	sub_wire118    <= data139x(39 DOWNTO 0);
	sub_wire117    <= data140x(39 DOWNTO 0);
	sub_wire116    <= data141x(39 DOWNTO 0);
	sub_wire115    <= data142x(39 DOWNTO 0);
	sub_wire114    <= data143x(39 DOWNTO 0);
	sub_wire113    <= data144x(39 DOWNTO 0);
	sub_wire112    <= data145x(39 DOWNTO 0);
	sub_wire111    <= data146x(39 DOWNTO 0);
	sub_wire110    <= data147x(39 DOWNTO 0);
	sub_wire109    <= data148x(39 DOWNTO 0);
	sub_wire108    <= data149x(39 DOWNTO 0);
	sub_wire107    <= data150x(39 DOWNTO 0);
	sub_wire106    <= data151x(39 DOWNTO 0);
	sub_wire105    <= data152x(39 DOWNTO 0);
	sub_wire104    <= data153x(39 DOWNTO 0);
	sub_wire103    <= data154x(39 DOWNTO 0);
	sub_wire102    <= data155x(39 DOWNTO 0);
	sub_wire101    <= data156x(39 DOWNTO 0);
	sub_wire100    <= data157x(39 DOWNTO 0);
	sub_wire99    <= data158x(39 DOWNTO 0);
	sub_wire98    <= data159x(39 DOWNTO 0);
	sub_wire97    <= data160x(39 DOWNTO 0);
	sub_wire96    <= data161x(39 DOWNTO 0);
	sub_wire95    <= data162x(39 DOWNTO 0);
	sub_wire94    <= data163x(39 DOWNTO 0);
	sub_wire93    <= data164x(39 DOWNTO 0);
	sub_wire92    <= data165x(39 DOWNTO 0);
	sub_wire91    <= data166x(39 DOWNTO 0);
	sub_wire90    <= data167x(39 DOWNTO 0);
	sub_wire89    <= data168x(39 DOWNTO 0);
	sub_wire88    <= data169x(39 DOWNTO 0);
	sub_wire87    <= data170x(39 DOWNTO 0);
	sub_wire86    <= data171x(39 DOWNTO 0);
	sub_wire85    <= data172x(39 DOWNTO 0);
	sub_wire84    <= data173x(39 DOWNTO 0);
	sub_wire83    <= data174x(39 DOWNTO 0);
	sub_wire82    <= data175x(39 DOWNTO 0);
	sub_wire81    <= data176x(39 DOWNTO 0);
	sub_wire80    <= data177x(39 DOWNTO 0);
	sub_wire79    <= data178x(39 DOWNTO 0);
	sub_wire78    <= data179x(39 DOWNTO 0);
	sub_wire77    <= data180x(39 DOWNTO 0);
	sub_wire76    <= data181x(39 DOWNTO 0);
	sub_wire75    <= data182x(39 DOWNTO 0);
	sub_wire74    <= data183x(39 DOWNTO 0);
	sub_wire73    <= data184x(39 DOWNTO 0);
	sub_wire72    <= data185x(39 DOWNTO 0);
	sub_wire71    <= data186x(39 DOWNTO 0);
	sub_wire70    <= data187x(39 DOWNTO 0);
	sub_wire69    <= data188x(39 DOWNTO 0);
	sub_wire68    <= data189x(39 DOWNTO 0);
	sub_wire67    <= data190x(39 DOWNTO 0);
	sub_wire66    <= data191x(39 DOWNTO 0);
	sub_wire65    <= data192x(39 DOWNTO 0);
	sub_wire64    <= data193x(39 DOWNTO 0);
	sub_wire63    <= data194x(39 DOWNTO 0);
	sub_wire62    <= data195x(39 DOWNTO 0);
	sub_wire61    <= data196x(39 DOWNTO 0);
	sub_wire60    <= data197x(39 DOWNTO 0);
	sub_wire59    <= data198x(39 DOWNTO 0);
	sub_wire58    <= data199x(39 DOWNTO 0);
	sub_wire57    <= data200x(39 DOWNTO 0);
	sub_wire56    <= data201x(39 DOWNTO 0);
	sub_wire55    <= data202x(39 DOWNTO 0);
	sub_wire54    <= data203x(39 DOWNTO 0);
	sub_wire53    <= data204x(39 DOWNTO 0);
	sub_wire52    <= data205x(39 DOWNTO 0);
	sub_wire51    <= data206x(39 DOWNTO 0);
	sub_wire50    <= data207x(39 DOWNTO 0);
	sub_wire49    <= data208x(39 DOWNTO 0);
	sub_wire48    <= data209x(39 DOWNTO 0);
	sub_wire47    <= data210x(39 DOWNTO 0);
	sub_wire46    <= data211x(39 DOWNTO 0);
	sub_wire45    <= data212x(39 DOWNTO 0);
	sub_wire44    <= data213x(39 DOWNTO 0);
	sub_wire43    <= data214x(39 DOWNTO 0);
	sub_wire42    <= data215x(39 DOWNTO 0);
	sub_wire41    <= data216x(39 DOWNTO 0);
	sub_wire40    <= data217x(39 DOWNTO 0);
	sub_wire39    <= data218x(39 DOWNTO 0);
	sub_wire38    <= data219x(39 DOWNTO 0);
	sub_wire37    <= data220x(39 DOWNTO 0);
	sub_wire36    <= data221x(39 DOWNTO 0);
	sub_wire35    <= data222x(39 DOWNTO 0);
	sub_wire34    <= data223x(39 DOWNTO 0);
	sub_wire33    <= data224x(39 DOWNTO 0);
	sub_wire32    <= data225x(39 DOWNTO 0);
	sub_wire31    <= data226x(39 DOWNTO 0);
	sub_wire30    <= data227x(39 DOWNTO 0);
	sub_wire29    <= data228x(39 DOWNTO 0);
	sub_wire28    <= data229x(39 DOWNTO 0);
	sub_wire27    <= data230x(39 DOWNTO 0);
	sub_wire26    <= data231x(39 DOWNTO 0);
	sub_wire25    <= data232x(39 DOWNTO 0);
	sub_wire24    <= data233x(39 DOWNTO 0);
	sub_wire23    <= data234x(39 DOWNTO 0);
	sub_wire22    <= data235x(39 DOWNTO 0);
	sub_wire21    <= data236x(39 DOWNTO 0);
	sub_wire20    <= data237x(39 DOWNTO 0);
	sub_wire19    <= data238x(39 DOWNTO 0);
	sub_wire18    <= data239x(39 DOWNTO 0);
	sub_wire17    <= data240x(39 DOWNTO 0);
	sub_wire16    <= data241x(39 DOWNTO 0);
	sub_wire15    <= data242x(39 DOWNTO 0);
	sub_wire14    <= data243x(39 DOWNTO 0);
	sub_wire13    <= data244x(39 DOWNTO 0);
	sub_wire12    <= data245x(39 DOWNTO 0);
	sub_wire11    <= data246x(39 DOWNTO 0);
	sub_wire10    <= data247x(39 DOWNTO 0);
	sub_wire9    <= data248x(39 DOWNTO 0);
	sub_wire8    <= data249x(39 DOWNTO 0);
	sub_wire7    <= data250x(39 DOWNTO 0);
	sub_wire6    <= data251x(39 DOWNTO 0);
	sub_wire5    <= data252x(39 DOWNTO 0);
	sub_wire4    <= data253x(39 DOWNTO 0);
	sub_wire3    <= data254x(39 DOWNTO 0);
	result    <= sub_wire0(39 DOWNTO 0);
	sub_wire1    <= data255x(39 DOWNTO 0);
	sub_wire2(255, 0)    <= sub_wire1(0);
	sub_wire2(255, 1)    <= sub_wire1(1);
	sub_wire2(255, 2)    <= sub_wire1(2);
	sub_wire2(255, 3)    <= sub_wire1(3);
	sub_wire2(255, 4)    <= sub_wire1(4);
	sub_wire2(255, 5)    <= sub_wire1(5);
	sub_wire2(255, 6)    <= sub_wire1(6);
	sub_wire2(255, 7)    <= sub_wire1(7);
	sub_wire2(255, 8)    <= sub_wire1(8);
	sub_wire2(255, 9)    <= sub_wire1(9);
	sub_wire2(255, 10)    <= sub_wire1(10);
	sub_wire2(255, 11)    <= sub_wire1(11);
	sub_wire2(255, 12)    <= sub_wire1(12);
	sub_wire2(255, 13)    <= sub_wire1(13);
	sub_wire2(255, 14)    <= sub_wire1(14);
	sub_wire2(255, 15)    <= sub_wire1(15);
	sub_wire2(255, 16)    <= sub_wire1(16);
	sub_wire2(255, 17)    <= sub_wire1(17);
	sub_wire2(255, 18)    <= sub_wire1(18);
	sub_wire2(255, 19)    <= sub_wire1(19);
	sub_wire2(255, 20)    <= sub_wire1(20);
	sub_wire2(255, 21)    <= sub_wire1(21);
	sub_wire2(255, 22)    <= sub_wire1(22);
	sub_wire2(255, 23)    <= sub_wire1(23);
	sub_wire2(255, 24)    <= sub_wire1(24);
	sub_wire2(255, 25)    <= sub_wire1(25);
	sub_wire2(255, 26)    <= sub_wire1(26);
	sub_wire2(255, 27)    <= sub_wire1(27);
	sub_wire2(255, 28)    <= sub_wire1(28);
	sub_wire2(255, 29)    <= sub_wire1(29);
	sub_wire2(255, 30)    <= sub_wire1(30);
	sub_wire2(255, 31)    <= sub_wire1(31);
	sub_wire2(255, 32)    <= sub_wire1(32);
	sub_wire2(255, 33)    <= sub_wire1(33);
	sub_wire2(255, 34)    <= sub_wire1(34);
	sub_wire2(255, 35)    <= sub_wire1(35);
	sub_wire2(255, 36)    <= sub_wire1(36);
	sub_wire2(255, 37)    <= sub_wire1(37);
	sub_wire2(255, 38)    <= sub_wire1(38);
	sub_wire2(255, 39)    <= sub_wire1(39);
	sub_wire2(254, 0)    <= sub_wire3(0);
	sub_wire2(254, 1)    <= sub_wire3(1);
	sub_wire2(254, 2)    <= sub_wire3(2);
	sub_wire2(254, 3)    <= sub_wire3(3);
	sub_wire2(254, 4)    <= sub_wire3(4);
	sub_wire2(254, 5)    <= sub_wire3(5);
	sub_wire2(254, 6)    <= sub_wire3(6);
	sub_wire2(254, 7)    <= sub_wire3(7);
	sub_wire2(254, 8)    <= sub_wire3(8);
	sub_wire2(254, 9)    <= sub_wire3(9);
	sub_wire2(254, 10)    <= sub_wire3(10);
	sub_wire2(254, 11)    <= sub_wire3(11);
	sub_wire2(254, 12)    <= sub_wire3(12);
	sub_wire2(254, 13)    <= sub_wire3(13);
	sub_wire2(254, 14)    <= sub_wire3(14);
	sub_wire2(254, 15)    <= sub_wire3(15);
	sub_wire2(254, 16)    <= sub_wire3(16);
	sub_wire2(254, 17)    <= sub_wire3(17);
	sub_wire2(254, 18)    <= sub_wire3(18);
	sub_wire2(254, 19)    <= sub_wire3(19);
	sub_wire2(254, 20)    <= sub_wire3(20);
	sub_wire2(254, 21)    <= sub_wire3(21);
	sub_wire2(254, 22)    <= sub_wire3(22);
	sub_wire2(254, 23)    <= sub_wire3(23);
	sub_wire2(254, 24)    <= sub_wire3(24);
	sub_wire2(254, 25)    <= sub_wire3(25);
	sub_wire2(254, 26)    <= sub_wire3(26);
	sub_wire2(254, 27)    <= sub_wire3(27);
	sub_wire2(254, 28)    <= sub_wire3(28);
	sub_wire2(254, 29)    <= sub_wire3(29);
	sub_wire2(254, 30)    <= sub_wire3(30);
	sub_wire2(254, 31)    <= sub_wire3(31);
	sub_wire2(254, 32)    <= sub_wire3(32);
	sub_wire2(254, 33)    <= sub_wire3(33);
	sub_wire2(254, 34)    <= sub_wire3(34);
	sub_wire2(254, 35)    <= sub_wire3(35);
	sub_wire2(254, 36)    <= sub_wire3(36);
	sub_wire2(254, 37)    <= sub_wire3(37);
	sub_wire2(254, 38)    <= sub_wire3(38);
	sub_wire2(254, 39)    <= sub_wire3(39);
	sub_wire2(253, 0)    <= sub_wire4(0);
	sub_wire2(253, 1)    <= sub_wire4(1);
	sub_wire2(253, 2)    <= sub_wire4(2);
	sub_wire2(253, 3)    <= sub_wire4(3);
	sub_wire2(253, 4)    <= sub_wire4(4);
	sub_wire2(253, 5)    <= sub_wire4(5);
	sub_wire2(253, 6)    <= sub_wire4(6);
	sub_wire2(253, 7)    <= sub_wire4(7);
	sub_wire2(253, 8)    <= sub_wire4(8);
	sub_wire2(253, 9)    <= sub_wire4(9);
	sub_wire2(253, 10)    <= sub_wire4(10);
	sub_wire2(253, 11)    <= sub_wire4(11);
	sub_wire2(253, 12)    <= sub_wire4(12);
	sub_wire2(253, 13)    <= sub_wire4(13);
	sub_wire2(253, 14)    <= sub_wire4(14);
	sub_wire2(253, 15)    <= sub_wire4(15);
	sub_wire2(253, 16)    <= sub_wire4(16);
	sub_wire2(253, 17)    <= sub_wire4(17);
	sub_wire2(253, 18)    <= sub_wire4(18);
	sub_wire2(253, 19)    <= sub_wire4(19);
	sub_wire2(253, 20)    <= sub_wire4(20);
	sub_wire2(253, 21)    <= sub_wire4(21);
	sub_wire2(253, 22)    <= sub_wire4(22);
	sub_wire2(253, 23)    <= sub_wire4(23);
	sub_wire2(253, 24)    <= sub_wire4(24);
	sub_wire2(253, 25)    <= sub_wire4(25);
	sub_wire2(253, 26)    <= sub_wire4(26);
	sub_wire2(253, 27)    <= sub_wire4(27);
	sub_wire2(253, 28)    <= sub_wire4(28);
	sub_wire2(253, 29)    <= sub_wire4(29);
	sub_wire2(253, 30)    <= sub_wire4(30);
	sub_wire2(253, 31)    <= sub_wire4(31);
	sub_wire2(253, 32)    <= sub_wire4(32);
	sub_wire2(253, 33)    <= sub_wire4(33);
	sub_wire2(253, 34)    <= sub_wire4(34);
	sub_wire2(253, 35)    <= sub_wire4(35);
	sub_wire2(253, 36)    <= sub_wire4(36);
	sub_wire2(253, 37)    <= sub_wire4(37);
	sub_wire2(253, 38)    <= sub_wire4(38);
	sub_wire2(253, 39)    <= sub_wire4(39);
	sub_wire2(252, 0)    <= sub_wire5(0);
	sub_wire2(252, 1)    <= sub_wire5(1);
	sub_wire2(252, 2)    <= sub_wire5(2);
	sub_wire2(252, 3)    <= sub_wire5(3);
	sub_wire2(252, 4)    <= sub_wire5(4);
	sub_wire2(252, 5)    <= sub_wire5(5);
	sub_wire2(252, 6)    <= sub_wire5(6);
	sub_wire2(252, 7)    <= sub_wire5(7);
	sub_wire2(252, 8)    <= sub_wire5(8);
	sub_wire2(252, 9)    <= sub_wire5(9);
	sub_wire2(252, 10)    <= sub_wire5(10);
	sub_wire2(252, 11)    <= sub_wire5(11);
	sub_wire2(252, 12)    <= sub_wire5(12);
	sub_wire2(252, 13)    <= sub_wire5(13);
	sub_wire2(252, 14)    <= sub_wire5(14);
	sub_wire2(252, 15)    <= sub_wire5(15);
	sub_wire2(252, 16)    <= sub_wire5(16);
	sub_wire2(252, 17)    <= sub_wire5(17);
	sub_wire2(252, 18)    <= sub_wire5(18);
	sub_wire2(252, 19)    <= sub_wire5(19);
	sub_wire2(252, 20)    <= sub_wire5(20);
	sub_wire2(252, 21)    <= sub_wire5(21);
	sub_wire2(252, 22)    <= sub_wire5(22);
	sub_wire2(252, 23)    <= sub_wire5(23);
	sub_wire2(252, 24)    <= sub_wire5(24);
	sub_wire2(252, 25)    <= sub_wire5(25);
	sub_wire2(252, 26)    <= sub_wire5(26);
	sub_wire2(252, 27)    <= sub_wire5(27);
	sub_wire2(252, 28)    <= sub_wire5(28);
	sub_wire2(252, 29)    <= sub_wire5(29);
	sub_wire2(252, 30)    <= sub_wire5(30);
	sub_wire2(252, 31)    <= sub_wire5(31);
	sub_wire2(252, 32)    <= sub_wire5(32);
	sub_wire2(252, 33)    <= sub_wire5(33);
	sub_wire2(252, 34)    <= sub_wire5(34);
	sub_wire2(252, 35)    <= sub_wire5(35);
	sub_wire2(252, 36)    <= sub_wire5(36);
	sub_wire2(252, 37)    <= sub_wire5(37);
	sub_wire2(252, 38)    <= sub_wire5(38);
	sub_wire2(252, 39)    <= sub_wire5(39);
	sub_wire2(251, 0)    <= sub_wire6(0);
	sub_wire2(251, 1)    <= sub_wire6(1);
	sub_wire2(251, 2)    <= sub_wire6(2);
	sub_wire2(251, 3)    <= sub_wire6(3);
	sub_wire2(251, 4)    <= sub_wire6(4);
	sub_wire2(251, 5)    <= sub_wire6(5);
	sub_wire2(251, 6)    <= sub_wire6(6);
	sub_wire2(251, 7)    <= sub_wire6(7);
	sub_wire2(251, 8)    <= sub_wire6(8);
	sub_wire2(251, 9)    <= sub_wire6(9);
	sub_wire2(251, 10)    <= sub_wire6(10);
	sub_wire2(251, 11)    <= sub_wire6(11);
	sub_wire2(251, 12)    <= sub_wire6(12);
	sub_wire2(251, 13)    <= sub_wire6(13);
	sub_wire2(251, 14)    <= sub_wire6(14);
	sub_wire2(251, 15)    <= sub_wire6(15);
	sub_wire2(251, 16)    <= sub_wire6(16);
	sub_wire2(251, 17)    <= sub_wire6(17);
	sub_wire2(251, 18)    <= sub_wire6(18);
	sub_wire2(251, 19)    <= sub_wire6(19);
	sub_wire2(251, 20)    <= sub_wire6(20);
	sub_wire2(251, 21)    <= sub_wire6(21);
	sub_wire2(251, 22)    <= sub_wire6(22);
	sub_wire2(251, 23)    <= sub_wire6(23);
	sub_wire2(251, 24)    <= sub_wire6(24);
	sub_wire2(251, 25)    <= sub_wire6(25);
	sub_wire2(251, 26)    <= sub_wire6(26);
	sub_wire2(251, 27)    <= sub_wire6(27);
	sub_wire2(251, 28)    <= sub_wire6(28);
	sub_wire2(251, 29)    <= sub_wire6(29);
	sub_wire2(251, 30)    <= sub_wire6(30);
	sub_wire2(251, 31)    <= sub_wire6(31);
	sub_wire2(251, 32)    <= sub_wire6(32);
	sub_wire2(251, 33)    <= sub_wire6(33);
	sub_wire2(251, 34)    <= sub_wire6(34);
	sub_wire2(251, 35)    <= sub_wire6(35);
	sub_wire2(251, 36)    <= sub_wire6(36);
	sub_wire2(251, 37)    <= sub_wire6(37);
	sub_wire2(251, 38)    <= sub_wire6(38);
	sub_wire2(251, 39)    <= sub_wire6(39);
	sub_wire2(250, 0)    <= sub_wire7(0);
	sub_wire2(250, 1)    <= sub_wire7(1);
	sub_wire2(250, 2)    <= sub_wire7(2);
	sub_wire2(250, 3)    <= sub_wire7(3);
	sub_wire2(250, 4)    <= sub_wire7(4);
	sub_wire2(250, 5)    <= sub_wire7(5);
	sub_wire2(250, 6)    <= sub_wire7(6);
	sub_wire2(250, 7)    <= sub_wire7(7);
	sub_wire2(250, 8)    <= sub_wire7(8);
	sub_wire2(250, 9)    <= sub_wire7(9);
	sub_wire2(250, 10)    <= sub_wire7(10);
	sub_wire2(250, 11)    <= sub_wire7(11);
	sub_wire2(250, 12)    <= sub_wire7(12);
	sub_wire2(250, 13)    <= sub_wire7(13);
	sub_wire2(250, 14)    <= sub_wire7(14);
	sub_wire2(250, 15)    <= sub_wire7(15);
	sub_wire2(250, 16)    <= sub_wire7(16);
	sub_wire2(250, 17)    <= sub_wire7(17);
	sub_wire2(250, 18)    <= sub_wire7(18);
	sub_wire2(250, 19)    <= sub_wire7(19);
	sub_wire2(250, 20)    <= sub_wire7(20);
	sub_wire2(250, 21)    <= sub_wire7(21);
	sub_wire2(250, 22)    <= sub_wire7(22);
	sub_wire2(250, 23)    <= sub_wire7(23);
	sub_wire2(250, 24)    <= sub_wire7(24);
	sub_wire2(250, 25)    <= sub_wire7(25);
	sub_wire2(250, 26)    <= sub_wire7(26);
	sub_wire2(250, 27)    <= sub_wire7(27);
	sub_wire2(250, 28)    <= sub_wire7(28);
	sub_wire2(250, 29)    <= sub_wire7(29);
	sub_wire2(250, 30)    <= sub_wire7(30);
	sub_wire2(250, 31)    <= sub_wire7(31);
	sub_wire2(250, 32)    <= sub_wire7(32);
	sub_wire2(250, 33)    <= sub_wire7(33);
	sub_wire2(250, 34)    <= sub_wire7(34);
	sub_wire2(250, 35)    <= sub_wire7(35);
	sub_wire2(250, 36)    <= sub_wire7(36);
	sub_wire2(250, 37)    <= sub_wire7(37);
	sub_wire2(250, 38)    <= sub_wire7(38);
	sub_wire2(250, 39)    <= sub_wire7(39);
	sub_wire2(249, 0)    <= sub_wire8(0);
	sub_wire2(249, 1)    <= sub_wire8(1);
	sub_wire2(249, 2)    <= sub_wire8(2);
	sub_wire2(249, 3)    <= sub_wire8(3);
	sub_wire2(249, 4)    <= sub_wire8(4);
	sub_wire2(249, 5)    <= sub_wire8(5);
	sub_wire2(249, 6)    <= sub_wire8(6);
	sub_wire2(249, 7)    <= sub_wire8(7);
	sub_wire2(249, 8)    <= sub_wire8(8);
	sub_wire2(249, 9)    <= sub_wire8(9);
	sub_wire2(249, 10)    <= sub_wire8(10);
	sub_wire2(249, 11)    <= sub_wire8(11);
	sub_wire2(249, 12)    <= sub_wire8(12);
	sub_wire2(249, 13)    <= sub_wire8(13);
	sub_wire2(249, 14)    <= sub_wire8(14);
	sub_wire2(249, 15)    <= sub_wire8(15);
	sub_wire2(249, 16)    <= sub_wire8(16);
	sub_wire2(249, 17)    <= sub_wire8(17);
	sub_wire2(249, 18)    <= sub_wire8(18);
	sub_wire2(249, 19)    <= sub_wire8(19);
	sub_wire2(249, 20)    <= sub_wire8(20);
	sub_wire2(249, 21)    <= sub_wire8(21);
	sub_wire2(249, 22)    <= sub_wire8(22);
	sub_wire2(249, 23)    <= sub_wire8(23);
	sub_wire2(249, 24)    <= sub_wire8(24);
	sub_wire2(249, 25)    <= sub_wire8(25);
	sub_wire2(249, 26)    <= sub_wire8(26);
	sub_wire2(249, 27)    <= sub_wire8(27);
	sub_wire2(249, 28)    <= sub_wire8(28);
	sub_wire2(249, 29)    <= sub_wire8(29);
	sub_wire2(249, 30)    <= sub_wire8(30);
	sub_wire2(249, 31)    <= sub_wire8(31);
	sub_wire2(249, 32)    <= sub_wire8(32);
	sub_wire2(249, 33)    <= sub_wire8(33);
	sub_wire2(249, 34)    <= sub_wire8(34);
	sub_wire2(249, 35)    <= sub_wire8(35);
	sub_wire2(249, 36)    <= sub_wire8(36);
	sub_wire2(249, 37)    <= sub_wire8(37);
	sub_wire2(249, 38)    <= sub_wire8(38);
	sub_wire2(249, 39)    <= sub_wire8(39);
	sub_wire2(248, 0)    <= sub_wire9(0);
	sub_wire2(248, 1)    <= sub_wire9(1);
	sub_wire2(248, 2)    <= sub_wire9(2);
	sub_wire2(248, 3)    <= sub_wire9(3);
	sub_wire2(248, 4)    <= sub_wire9(4);
	sub_wire2(248, 5)    <= sub_wire9(5);
	sub_wire2(248, 6)    <= sub_wire9(6);
	sub_wire2(248, 7)    <= sub_wire9(7);
	sub_wire2(248, 8)    <= sub_wire9(8);
	sub_wire2(248, 9)    <= sub_wire9(9);
	sub_wire2(248, 10)    <= sub_wire9(10);
	sub_wire2(248, 11)    <= sub_wire9(11);
	sub_wire2(248, 12)    <= sub_wire9(12);
	sub_wire2(248, 13)    <= sub_wire9(13);
	sub_wire2(248, 14)    <= sub_wire9(14);
	sub_wire2(248, 15)    <= sub_wire9(15);
	sub_wire2(248, 16)    <= sub_wire9(16);
	sub_wire2(248, 17)    <= sub_wire9(17);
	sub_wire2(248, 18)    <= sub_wire9(18);
	sub_wire2(248, 19)    <= sub_wire9(19);
	sub_wire2(248, 20)    <= sub_wire9(20);
	sub_wire2(248, 21)    <= sub_wire9(21);
	sub_wire2(248, 22)    <= sub_wire9(22);
	sub_wire2(248, 23)    <= sub_wire9(23);
	sub_wire2(248, 24)    <= sub_wire9(24);
	sub_wire2(248, 25)    <= sub_wire9(25);
	sub_wire2(248, 26)    <= sub_wire9(26);
	sub_wire2(248, 27)    <= sub_wire9(27);
	sub_wire2(248, 28)    <= sub_wire9(28);
	sub_wire2(248, 29)    <= sub_wire9(29);
	sub_wire2(248, 30)    <= sub_wire9(30);
	sub_wire2(248, 31)    <= sub_wire9(31);
	sub_wire2(248, 32)    <= sub_wire9(32);
	sub_wire2(248, 33)    <= sub_wire9(33);
	sub_wire2(248, 34)    <= sub_wire9(34);
	sub_wire2(248, 35)    <= sub_wire9(35);
	sub_wire2(248, 36)    <= sub_wire9(36);
	sub_wire2(248, 37)    <= sub_wire9(37);
	sub_wire2(248, 38)    <= sub_wire9(38);
	sub_wire2(248, 39)    <= sub_wire9(39);
	sub_wire2(247, 0)    <= sub_wire10(0);
	sub_wire2(247, 1)    <= sub_wire10(1);
	sub_wire2(247, 2)    <= sub_wire10(2);
	sub_wire2(247, 3)    <= sub_wire10(3);
	sub_wire2(247, 4)    <= sub_wire10(4);
	sub_wire2(247, 5)    <= sub_wire10(5);
	sub_wire2(247, 6)    <= sub_wire10(6);
	sub_wire2(247, 7)    <= sub_wire10(7);
	sub_wire2(247, 8)    <= sub_wire10(8);
	sub_wire2(247, 9)    <= sub_wire10(9);
	sub_wire2(247, 10)    <= sub_wire10(10);
	sub_wire2(247, 11)    <= sub_wire10(11);
	sub_wire2(247, 12)    <= sub_wire10(12);
	sub_wire2(247, 13)    <= sub_wire10(13);
	sub_wire2(247, 14)    <= sub_wire10(14);
	sub_wire2(247, 15)    <= sub_wire10(15);
	sub_wire2(247, 16)    <= sub_wire10(16);
	sub_wire2(247, 17)    <= sub_wire10(17);
	sub_wire2(247, 18)    <= sub_wire10(18);
	sub_wire2(247, 19)    <= sub_wire10(19);
	sub_wire2(247, 20)    <= sub_wire10(20);
	sub_wire2(247, 21)    <= sub_wire10(21);
	sub_wire2(247, 22)    <= sub_wire10(22);
	sub_wire2(247, 23)    <= sub_wire10(23);
	sub_wire2(247, 24)    <= sub_wire10(24);
	sub_wire2(247, 25)    <= sub_wire10(25);
	sub_wire2(247, 26)    <= sub_wire10(26);
	sub_wire2(247, 27)    <= sub_wire10(27);
	sub_wire2(247, 28)    <= sub_wire10(28);
	sub_wire2(247, 29)    <= sub_wire10(29);
	sub_wire2(247, 30)    <= sub_wire10(30);
	sub_wire2(247, 31)    <= sub_wire10(31);
	sub_wire2(247, 32)    <= sub_wire10(32);
	sub_wire2(247, 33)    <= sub_wire10(33);
	sub_wire2(247, 34)    <= sub_wire10(34);
	sub_wire2(247, 35)    <= sub_wire10(35);
	sub_wire2(247, 36)    <= sub_wire10(36);
	sub_wire2(247, 37)    <= sub_wire10(37);
	sub_wire2(247, 38)    <= sub_wire10(38);
	sub_wire2(247, 39)    <= sub_wire10(39);
	sub_wire2(246, 0)    <= sub_wire11(0);
	sub_wire2(246, 1)    <= sub_wire11(1);
	sub_wire2(246, 2)    <= sub_wire11(2);
	sub_wire2(246, 3)    <= sub_wire11(3);
	sub_wire2(246, 4)    <= sub_wire11(4);
	sub_wire2(246, 5)    <= sub_wire11(5);
	sub_wire2(246, 6)    <= sub_wire11(6);
	sub_wire2(246, 7)    <= sub_wire11(7);
	sub_wire2(246, 8)    <= sub_wire11(8);
	sub_wire2(246, 9)    <= sub_wire11(9);
	sub_wire2(246, 10)    <= sub_wire11(10);
	sub_wire2(246, 11)    <= sub_wire11(11);
	sub_wire2(246, 12)    <= sub_wire11(12);
	sub_wire2(246, 13)    <= sub_wire11(13);
	sub_wire2(246, 14)    <= sub_wire11(14);
	sub_wire2(246, 15)    <= sub_wire11(15);
	sub_wire2(246, 16)    <= sub_wire11(16);
	sub_wire2(246, 17)    <= sub_wire11(17);
	sub_wire2(246, 18)    <= sub_wire11(18);
	sub_wire2(246, 19)    <= sub_wire11(19);
	sub_wire2(246, 20)    <= sub_wire11(20);
	sub_wire2(246, 21)    <= sub_wire11(21);
	sub_wire2(246, 22)    <= sub_wire11(22);
	sub_wire2(246, 23)    <= sub_wire11(23);
	sub_wire2(246, 24)    <= sub_wire11(24);
	sub_wire2(246, 25)    <= sub_wire11(25);
	sub_wire2(246, 26)    <= sub_wire11(26);
	sub_wire2(246, 27)    <= sub_wire11(27);
	sub_wire2(246, 28)    <= sub_wire11(28);
	sub_wire2(246, 29)    <= sub_wire11(29);
	sub_wire2(246, 30)    <= sub_wire11(30);
	sub_wire2(246, 31)    <= sub_wire11(31);
	sub_wire2(246, 32)    <= sub_wire11(32);
	sub_wire2(246, 33)    <= sub_wire11(33);
	sub_wire2(246, 34)    <= sub_wire11(34);
	sub_wire2(246, 35)    <= sub_wire11(35);
	sub_wire2(246, 36)    <= sub_wire11(36);
	sub_wire2(246, 37)    <= sub_wire11(37);
	sub_wire2(246, 38)    <= sub_wire11(38);
	sub_wire2(246, 39)    <= sub_wire11(39);
	sub_wire2(245, 0)    <= sub_wire12(0);
	sub_wire2(245, 1)    <= sub_wire12(1);
	sub_wire2(245, 2)    <= sub_wire12(2);
	sub_wire2(245, 3)    <= sub_wire12(3);
	sub_wire2(245, 4)    <= sub_wire12(4);
	sub_wire2(245, 5)    <= sub_wire12(5);
	sub_wire2(245, 6)    <= sub_wire12(6);
	sub_wire2(245, 7)    <= sub_wire12(7);
	sub_wire2(245, 8)    <= sub_wire12(8);
	sub_wire2(245, 9)    <= sub_wire12(9);
	sub_wire2(245, 10)    <= sub_wire12(10);
	sub_wire2(245, 11)    <= sub_wire12(11);
	sub_wire2(245, 12)    <= sub_wire12(12);
	sub_wire2(245, 13)    <= sub_wire12(13);
	sub_wire2(245, 14)    <= sub_wire12(14);
	sub_wire2(245, 15)    <= sub_wire12(15);
	sub_wire2(245, 16)    <= sub_wire12(16);
	sub_wire2(245, 17)    <= sub_wire12(17);
	sub_wire2(245, 18)    <= sub_wire12(18);
	sub_wire2(245, 19)    <= sub_wire12(19);
	sub_wire2(245, 20)    <= sub_wire12(20);
	sub_wire2(245, 21)    <= sub_wire12(21);
	sub_wire2(245, 22)    <= sub_wire12(22);
	sub_wire2(245, 23)    <= sub_wire12(23);
	sub_wire2(245, 24)    <= sub_wire12(24);
	sub_wire2(245, 25)    <= sub_wire12(25);
	sub_wire2(245, 26)    <= sub_wire12(26);
	sub_wire2(245, 27)    <= sub_wire12(27);
	sub_wire2(245, 28)    <= sub_wire12(28);
	sub_wire2(245, 29)    <= sub_wire12(29);
	sub_wire2(245, 30)    <= sub_wire12(30);
	sub_wire2(245, 31)    <= sub_wire12(31);
	sub_wire2(245, 32)    <= sub_wire12(32);
	sub_wire2(245, 33)    <= sub_wire12(33);
	sub_wire2(245, 34)    <= sub_wire12(34);
	sub_wire2(245, 35)    <= sub_wire12(35);
	sub_wire2(245, 36)    <= sub_wire12(36);
	sub_wire2(245, 37)    <= sub_wire12(37);
	sub_wire2(245, 38)    <= sub_wire12(38);
	sub_wire2(245, 39)    <= sub_wire12(39);
	sub_wire2(244, 0)    <= sub_wire13(0);
	sub_wire2(244, 1)    <= sub_wire13(1);
	sub_wire2(244, 2)    <= sub_wire13(2);
	sub_wire2(244, 3)    <= sub_wire13(3);
	sub_wire2(244, 4)    <= sub_wire13(4);
	sub_wire2(244, 5)    <= sub_wire13(5);
	sub_wire2(244, 6)    <= sub_wire13(6);
	sub_wire2(244, 7)    <= sub_wire13(7);
	sub_wire2(244, 8)    <= sub_wire13(8);
	sub_wire2(244, 9)    <= sub_wire13(9);
	sub_wire2(244, 10)    <= sub_wire13(10);
	sub_wire2(244, 11)    <= sub_wire13(11);
	sub_wire2(244, 12)    <= sub_wire13(12);
	sub_wire2(244, 13)    <= sub_wire13(13);
	sub_wire2(244, 14)    <= sub_wire13(14);
	sub_wire2(244, 15)    <= sub_wire13(15);
	sub_wire2(244, 16)    <= sub_wire13(16);
	sub_wire2(244, 17)    <= sub_wire13(17);
	sub_wire2(244, 18)    <= sub_wire13(18);
	sub_wire2(244, 19)    <= sub_wire13(19);
	sub_wire2(244, 20)    <= sub_wire13(20);
	sub_wire2(244, 21)    <= sub_wire13(21);
	sub_wire2(244, 22)    <= sub_wire13(22);
	sub_wire2(244, 23)    <= sub_wire13(23);
	sub_wire2(244, 24)    <= sub_wire13(24);
	sub_wire2(244, 25)    <= sub_wire13(25);
	sub_wire2(244, 26)    <= sub_wire13(26);
	sub_wire2(244, 27)    <= sub_wire13(27);
	sub_wire2(244, 28)    <= sub_wire13(28);
	sub_wire2(244, 29)    <= sub_wire13(29);
	sub_wire2(244, 30)    <= sub_wire13(30);
	sub_wire2(244, 31)    <= sub_wire13(31);
	sub_wire2(244, 32)    <= sub_wire13(32);
	sub_wire2(244, 33)    <= sub_wire13(33);
	sub_wire2(244, 34)    <= sub_wire13(34);
	sub_wire2(244, 35)    <= sub_wire13(35);
	sub_wire2(244, 36)    <= sub_wire13(36);
	sub_wire2(244, 37)    <= sub_wire13(37);
	sub_wire2(244, 38)    <= sub_wire13(38);
	sub_wire2(244, 39)    <= sub_wire13(39);
	sub_wire2(243, 0)    <= sub_wire14(0);
	sub_wire2(243, 1)    <= sub_wire14(1);
	sub_wire2(243, 2)    <= sub_wire14(2);
	sub_wire2(243, 3)    <= sub_wire14(3);
	sub_wire2(243, 4)    <= sub_wire14(4);
	sub_wire2(243, 5)    <= sub_wire14(5);
	sub_wire2(243, 6)    <= sub_wire14(6);
	sub_wire2(243, 7)    <= sub_wire14(7);
	sub_wire2(243, 8)    <= sub_wire14(8);
	sub_wire2(243, 9)    <= sub_wire14(9);
	sub_wire2(243, 10)    <= sub_wire14(10);
	sub_wire2(243, 11)    <= sub_wire14(11);
	sub_wire2(243, 12)    <= sub_wire14(12);
	sub_wire2(243, 13)    <= sub_wire14(13);
	sub_wire2(243, 14)    <= sub_wire14(14);
	sub_wire2(243, 15)    <= sub_wire14(15);
	sub_wire2(243, 16)    <= sub_wire14(16);
	sub_wire2(243, 17)    <= sub_wire14(17);
	sub_wire2(243, 18)    <= sub_wire14(18);
	sub_wire2(243, 19)    <= sub_wire14(19);
	sub_wire2(243, 20)    <= sub_wire14(20);
	sub_wire2(243, 21)    <= sub_wire14(21);
	sub_wire2(243, 22)    <= sub_wire14(22);
	sub_wire2(243, 23)    <= sub_wire14(23);
	sub_wire2(243, 24)    <= sub_wire14(24);
	sub_wire2(243, 25)    <= sub_wire14(25);
	sub_wire2(243, 26)    <= sub_wire14(26);
	sub_wire2(243, 27)    <= sub_wire14(27);
	sub_wire2(243, 28)    <= sub_wire14(28);
	sub_wire2(243, 29)    <= sub_wire14(29);
	sub_wire2(243, 30)    <= sub_wire14(30);
	sub_wire2(243, 31)    <= sub_wire14(31);
	sub_wire2(243, 32)    <= sub_wire14(32);
	sub_wire2(243, 33)    <= sub_wire14(33);
	sub_wire2(243, 34)    <= sub_wire14(34);
	sub_wire2(243, 35)    <= sub_wire14(35);
	sub_wire2(243, 36)    <= sub_wire14(36);
	sub_wire2(243, 37)    <= sub_wire14(37);
	sub_wire2(243, 38)    <= sub_wire14(38);
	sub_wire2(243, 39)    <= sub_wire14(39);
	sub_wire2(242, 0)    <= sub_wire15(0);
	sub_wire2(242, 1)    <= sub_wire15(1);
	sub_wire2(242, 2)    <= sub_wire15(2);
	sub_wire2(242, 3)    <= sub_wire15(3);
	sub_wire2(242, 4)    <= sub_wire15(4);
	sub_wire2(242, 5)    <= sub_wire15(5);
	sub_wire2(242, 6)    <= sub_wire15(6);
	sub_wire2(242, 7)    <= sub_wire15(7);
	sub_wire2(242, 8)    <= sub_wire15(8);
	sub_wire2(242, 9)    <= sub_wire15(9);
	sub_wire2(242, 10)    <= sub_wire15(10);
	sub_wire2(242, 11)    <= sub_wire15(11);
	sub_wire2(242, 12)    <= sub_wire15(12);
	sub_wire2(242, 13)    <= sub_wire15(13);
	sub_wire2(242, 14)    <= sub_wire15(14);
	sub_wire2(242, 15)    <= sub_wire15(15);
	sub_wire2(242, 16)    <= sub_wire15(16);
	sub_wire2(242, 17)    <= sub_wire15(17);
	sub_wire2(242, 18)    <= sub_wire15(18);
	sub_wire2(242, 19)    <= sub_wire15(19);
	sub_wire2(242, 20)    <= sub_wire15(20);
	sub_wire2(242, 21)    <= sub_wire15(21);
	sub_wire2(242, 22)    <= sub_wire15(22);
	sub_wire2(242, 23)    <= sub_wire15(23);
	sub_wire2(242, 24)    <= sub_wire15(24);
	sub_wire2(242, 25)    <= sub_wire15(25);
	sub_wire2(242, 26)    <= sub_wire15(26);
	sub_wire2(242, 27)    <= sub_wire15(27);
	sub_wire2(242, 28)    <= sub_wire15(28);
	sub_wire2(242, 29)    <= sub_wire15(29);
	sub_wire2(242, 30)    <= sub_wire15(30);
	sub_wire2(242, 31)    <= sub_wire15(31);
	sub_wire2(242, 32)    <= sub_wire15(32);
	sub_wire2(242, 33)    <= sub_wire15(33);
	sub_wire2(242, 34)    <= sub_wire15(34);
	sub_wire2(242, 35)    <= sub_wire15(35);
	sub_wire2(242, 36)    <= sub_wire15(36);
	sub_wire2(242, 37)    <= sub_wire15(37);
	sub_wire2(242, 38)    <= sub_wire15(38);
	sub_wire2(242, 39)    <= sub_wire15(39);
	sub_wire2(241, 0)    <= sub_wire16(0);
	sub_wire2(241, 1)    <= sub_wire16(1);
	sub_wire2(241, 2)    <= sub_wire16(2);
	sub_wire2(241, 3)    <= sub_wire16(3);
	sub_wire2(241, 4)    <= sub_wire16(4);
	sub_wire2(241, 5)    <= sub_wire16(5);
	sub_wire2(241, 6)    <= sub_wire16(6);
	sub_wire2(241, 7)    <= sub_wire16(7);
	sub_wire2(241, 8)    <= sub_wire16(8);
	sub_wire2(241, 9)    <= sub_wire16(9);
	sub_wire2(241, 10)    <= sub_wire16(10);
	sub_wire2(241, 11)    <= sub_wire16(11);
	sub_wire2(241, 12)    <= sub_wire16(12);
	sub_wire2(241, 13)    <= sub_wire16(13);
	sub_wire2(241, 14)    <= sub_wire16(14);
	sub_wire2(241, 15)    <= sub_wire16(15);
	sub_wire2(241, 16)    <= sub_wire16(16);
	sub_wire2(241, 17)    <= sub_wire16(17);
	sub_wire2(241, 18)    <= sub_wire16(18);
	sub_wire2(241, 19)    <= sub_wire16(19);
	sub_wire2(241, 20)    <= sub_wire16(20);
	sub_wire2(241, 21)    <= sub_wire16(21);
	sub_wire2(241, 22)    <= sub_wire16(22);
	sub_wire2(241, 23)    <= sub_wire16(23);
	sub_wire2(241, 24)    <= sub_wire16(24);
	sub_wire2(241, 25)    <= sub_wire16(25);
	sub_wire2(241, 26)    <= sub_wire16(26);
	sub_wire2(241, 27)    <= sub_wire16(27);
	sub_wire2(241, 28)    <= sub_wire16(28);
	sub_wire2(241, 29)    <= sub_wire16(29);
	sub_wire2(241, 30)    <= sub_wire16(30);
	sub_wire2(241, 31)    <= sub_wire16(31);
	sub_wire2(241, 32)    <= sub_wire16(32);
	sub_wire2(241, 33)    <= sub_wire16(33);
	sub_wire2(241, 34)    <= sub_wire16(34);
	sub_wire2(241, 35)    <= sub_wire16(35);
	sub_wire2(241, 36)    <= sub_wire16(36);
	sub_wire2(241, 37)    <= sub_wire16(37);
	sub_wire2(241, 38)    <= sub_wire16(38);
	sub_wire2(241, 39)    <= sub_wire16(39);
	sub_wire2(240, 0)    <= sub_wire17(0);
	sub_wire2(240, 1)    <= sub_wire17(1);
	sub_wire2(240, 2)    <= sub_wire17(2);
	sub_wire2(240, 3)    <= sub_wire17(3);
	sub_wire2(240, 4)    <= sub_wire17(4);
	sub_wire2(240, 5)    <= sub_wire17(5);
	sub_wire2(240, 6)    <= sub_wire17(6);
	sub_wire2(240, 7)    <= sub_wire17(7);
	sub_wire2(240, 8)    <= sub_wire17(8);
	sub_wire2(240, 9)    <= sub_wire17(9);
	sub_wire2(240, 10)    <= sub_wire17(10);
	sub_wire2(240, 11)    <= sub_wire17(11);
	sub_wire2(240, 12)    <= sub_wire17(12);
	sub_wire2(240, 13)    <= sub_wire17(13);
	sub_wire2(240, 14)    <= sub_wire17(14);
	sub_wire2(240, 15)    <= sub_wire17(15);
	sub_wire2(240, 16)    <= sub_wire17(16);
	sub_wire2(240, 17)    <= sub_wire17(17);
	sub_wire2(240, 18)    <= sub_wire17(18);
	sub_wire2(240, 19)    <= sub_wire17(19);
	sub_wire2(240, 20)    <= sub_wire17(20);
	sub_wire2(240, 21)    <= sub_wire17(21);
	sub_wire2(240, 22)    <= sub_wire17(22);
	sub_wire2(240, 23)    <= sub_wire17(23);
	sub_wire2(240, 24)    <= sub_wire17(24);
	sub_wire2(240, 25)    <= sub_wire17(25);
	sub_wire2(240, 26)    <= sub_wire17(26);
	sub_wire2(240, 27)    <= sub_wire17(27);
	sub_wire2(240, 28)    <= sub_wire17(28);
	sub_wire2(240, 29)    <= sub_wire17(29);
	sub_wire2(240, 30)    <= sub_wire17(30);
	sub_wire2(240, 31)    <= sub_wire17(31);
	sub_wire2(240, 32)    <= sub_wire17(32);
	sub_wire2(240, 33)    <= sub_wire17(33);
	sub_wire2(240, 34)    <= sub_wire17(34);
	sub_wire2(240, 35)    <= sub_wire17(35);
	sub_wire2(240, 36)    <= sub_wire17(36);
	sub_wire2(240, 37)    <= sub_wire17(37);
	sub_wire2(240, 38)    <= sub_wire17(38);
	sub_wire2(240, 39)    <= sub_wire17(39);
	sub_wire2(239, 0)    <= sub_wire18(0);
	sub_wire2(239, 1)    <= sub_wire18(1);
	sub_wire2(239, 2)    <= sub_wire18(2);
	sub_wire2(239, 3)    <= sub_wire18(3);
	sub_wire2(239, 4)    <= sub_wire18(4);
	sub_wire2(239, 5)    <= sub_wire18(5);
	sub_wire2(239, 6)    <= sub_wire18(6);
	sub_wire2(239, 7)    <= sub_wire18(7);
	sub_wire2(239, 8)    <= sub_wire18(8);
	sub_wire2(239, 9)    <= sub_wire18(9);
	sub_wire2(239, 10)    <= sub_wire18(10);
	sub_wire2(239, 11)    <= sub_wire18(11);
	sub_wire2(239, 12)    <= sub_wire18(12);
	sub_wire2(239, 13)    <= sub_wire18(13);
	sub_wire2(239, 14)    <= sub_wire18(14);
	sub_wire2(239, 15)    <= sub_wire18(15);
	sub_wire2(239, 16)    <= sub_wire18(16);
	sub_wire2(239, 17)    <= sub_wire18(17);
	sub_wire2(239, 18)    <= sub_wire18(18);
	sub_wire2(239, 19)    <= sub_wire18(19);
	sub_wire2(239, 20)    <= sub_wire18(20);
	sub_wire2(239, 21)    <= sub_wire18(21);
	sub_wire2(239, 22)    <= sub_wire18(22);
	sub_wire2(239, 23)    <= sub_wire18(23);
	sub_wire2(239, 24)    <= sub_wire18(24);
	sub_wire2(239, 25)    <= sub_wire18(25);
	sub_wire2(239, 26)    <= sub_wire18(26);
	sub_wire2(239, 27)    <= sub_wire18(27);
	sub_wire2(239, 28)    <= sub_wire18(28);
	sub_wire2(239, 29)    <= sub_wire18(29);
	sub_wire2(239, 30)    <= sub_wire18(30);
	sub_wire2(239, 31)    <= sub_wire18(31);
	sub_wire2(239, 32)    <= sub_wire18(32);
	sub_wire2(239, 33)    <= sub_wire18(33);
	sub_wire2(239, 34)    <= sub_wire18(34);
	sub_wire2(239, 35)    <= sub_wire18(35);
	sub_wire2(239, 36)    <= sub_wire18(36);
	sub_wire2(239, 37)    <= sub_wire18(37);
	sub_wire2(239, 38)    <= sub_wire18(38);
	sub_wire2(239, 39)    <= sub_wire18(39);
	sub_wire2(238, 0)    <= sub_wire19(0);
	sub_wire2(238, 1)    <= sub_wire19(1);
	sub_wire2(238, 2)    <= sub_wire19(2);
	sub_wire2(238, 3)    <= sub_wire19(3);
	sub_wire2(238, 4)    <= sub_wire19(4);
	sub_wire2(238, 5)    <= sub_wire19(5);
	sub_wire2(238, 6)    <= sub_wire19(6);
	sub_wire2(238, 7)    <= sub_wire19(7);
	sub_wire2(238, 8)    <= sub_wire19(8);
	sub_wire2(238, 9)    <= sub_wire19(9);
	sub_wire2(238, 10)    <= sub_wire19(10);
	sub_wire2(238, 11)    <= sub_wire19(11);
	sub_wire2(238, 12)    <= sub_wire19(12);
	sub_wire2(238, 13)    <= sub_wire19(13);
	sub_wire2(238, 14)    <= sub_wire19(14);
	sub_wire2(238, 15)    <= sub_wire19(15);
	sub_wire2(238, 16)    <= sub_wire19(16);
	sub_wire2(238, 17)    <= sub_wire19(17);
	sub_wire2(238, 18)    <= sub_wire19(18);
	sub_wire2(238, 19)    <= sub_wire19(19);
	sub_wire2(238, 20)    <= sub_wire19(20);
	sub_wire2(238, 21)    <= sub_wire19(21);
	sub_wire2(238, 22)    <= sub_wire19(22);
	sub_wire2(238, 23)    <= sub_wire19(23);
	sub_wire2(238, 24)    <= sub_wire19(24);
	sub_wire2(238, 25)    <= sub_wire19(25);
	sub_wire2(238, 26)    <= sub_wire19(26);
	sub_wire2(238, 27)    <= sub_wire19(27);
	sub_wire2(238, 28)    <= sub_wire19(28);
	sub_wire2(238, 29)    <= sub_wire19(29);
	sub_wire2(238, 30)    <= sub_wire19(30);
	sub_wire2(238, 31)    <= sub_wire19(31);
	sub_wire2(238, 32)    <= sub_wire19(32);
	sub_wire2(238, 33)    <= sub_wire19(33);
	sub_wire2(238, 34)    <= sub_wire19(34);
	sub_wire2(238, 35)    <= sub_wire19(35);
	sub_wire2(238, 36)    <= sub_wire19(36);
	sub_wire2(238, 37)    <= sub_wire19(37);
	sub_wire2(238, 38)    <= sub_wire19(38);
	sub_wire2(238, 39)    <= sub_wire19(39);
	sub_wire2(237, 0)    <= sub_wire20(0);
	sub_wire2(237, 1)    <= sub_wire20(1);
	sub_wire2(237, 2)    <= sub_wire20(2);
	sub_wire2(237, 3)    <= sub_wire20(3);
	sub_wire2(237, 4)    <= sub_wire20(4);
	sub_wire2(237, 5)    <= sub_wire20(5);
	sub_wire2(237, 6)    <= sub_wire20(6);
	sub_wire2(237, 7)    <= sub_wire20(7);
	sub_wire2(237, 8)    <= sub_wire20(8);
	sub_wire2(237, 9)    <= sub_wire20(9);
	sub_wire2(237, 10)    <= sub_wire20(10);
	sub_wire2(237, 11)    <= sub_wire20(11);
	sub_wire2(237, 12)    <= sub_wire20(12);
	sub_wire2(237, 13)    <= sub_wire20(13);
	sub_wire2(237, 14)    <= sub_wire20(14);
	sub_wire2(237, 15)    <= sub_wire20(15);
	sub_wire2(237, 16)    <= sub_wire20(16);
	sub_wire2(237, 17)    <= sub_wire20(17);
	sub_wire2(237, 18)    <= sub_wire20(18);
	sub_wire2(237, 19)    <= sub_wire20(19);
	sub_wire2(237, 20)    <= sub_wire20(20);
	sub_wire2(237, 21)    <= sub_wire20(21);
	sub_wire2(237, 22)    <= sub_wire20(22);
	sub_wire2(237, 23)    <= sub_wire20(23);
	sub_wire2(237, 24)    <= sub_wire20(24);
	sub_wire2(237, 25)    <= sub_wire20(25);
	sub_wire2(237, 26)    <= sub_wire20(26);
	sub_wire2(237, 27)    <= sub_wire20(27);
	sub_wire2(237, 28)    <= sub_wire20(28);
	sub_wire2(237, 29)    <= sub_wire20(29);
	sub_wire2(237, 30)    <= sub_wire20(30);
	sub_wire2(237, 31)    <= sub_wire20(31);
	sub_wire2(237, 32)    <= sub_wire20(32);
	sub_wire2(237, 33)    <= sub_wire20(33);
	sub_wire2(237, 34)    <= sub_wire20(34);
	sub_wire2(237, 35)    <= sub_wire20(35);
	sub_wire2(237, 36)    <= sub_wire20(36);
	sub_wire2(237, 37)    <= sub_wire20(37);
	sub_wire2(237, 38)    <= sub_wire20(38);
	sub_wire2(237, 39)    <= sub_wire20(39);
	sub_wire2(236, 0)    <= sub_wire21(0);
	sub_wire2(236, 1)    <= sub_wire21(1);
	sub_wire2(236, 2)    <= sub_wire21(2);
	sub_wire2(236, 3)    <= sub_wire21(3);
	sub_wire2(236, 4)    <= sub_wire21(4);
	sub_wire2(236, 5)    <= sub_wire21(5);
	sub_wire2(236, 6)    <= sub_wire21(6);
	sub_wire2(236, 7)    <= sub_wire21(7);
	sub_wire2(236, 8)    <= sub_wire21(8);
	sub_wire2(236, 9)    <= sub_wire21(9);
	sub_wire2(236, 10)    <= sub_wire21(10);
	sub_wire2(236, 11)    <= sub_wire21(11);
	sub_wire2(236, 12)    <= sub_wire21(12);
	sub_wire2(236, 13)    <= sub_wire21(13);
	sub_wire2(236, 14)    <= sub_wire21(14);
	sub_wire2(236, 15)    <= sub_wire21(15);
	sub_wire2(236, 16)    <= sub_wire21(16);
	sub_wire2(236, 17)    <= sub_wire21(17);
	sub_wire2(236, 18)    <= sub_wire21(18);
	sub_wire2(236, 19)    <= sub_wire21(19);
	sub_wire2(236, 20)    <= sub_wire21(20);
	sub_wire2(236, 21)    <= sub_wire21(21);
	sub_wire2(236, 22)    <= sub_wire21(22);
	sub_wire2(236, 23)    <= sub_wire21(23);
	sub_wire2(236, 24)    <= sub_wire21(24);
	sub_wire2(236, 25)    <= sub_wire21(25);
	sub_wire2(236, 26)    <= sub_wire21(26);
	sub_wire2(236, 27)    <= sub_wire21(27);
	sub_wire2(236, 28)    <= sub_wire21(28);
	sub_wire2(236, 29)    <= sub_wire21(29);
	sub_wire2(236, 30)    <= sub_wire21(30);
	sub_wire2(236, 31)    <= sub_wire21(31);
	sub_wire2(236, 32)    <= sub_wire21(32);
	sub_wire2(236, 33)    <= sub_wire21(33);
	sub_wire2(236, 34)    <= sub_wire21(34);
	sub_wire2(236, 35)    <= sub_wire21(35);
	sub_wire2(236, 36)    <= sub_wire21(36);
	sub_wire2(236, 37)    <= sub_wire21(37);
	sub_wire2(236, 38)    <= sub_wire21(38);
	sub_wire2(236, 39)    <= sub_wire21(39);
	sub_wire2(235, 0)    <= sub_wire22(0);
	sub_wire2(235, 1)    <= sub_wire22(1);
	sub_wire2(235, 2)    <= sub_wire22(2);
	sub_wire2(235, 3)    <= sub_wire22(3);
	sub_wire2(235, 4)    <= sub_wire22(4);
	sub_wire2(235, 5)    <= sub_wire22(5);
	sub_wire2(235, 6)    <= sub_wire22(6);
	sub_wire2(235, 7)    <= sub_wire22(7);
	sub_wire2(235, 8)    <= sub_wire22(8);
	sub_wire2(235, 9)    <= sub_wire22(9);
	sub_wire2(235, 10)    <= sub_wire22(10);
	sub_wire2(235, 11)    <= sub_wire22(11);
	sub_wire2(235, 12)    <= sub_wire22(12);
	sub_wire2(235, 13)    <= sub_wire22(13);
	sub_wire2(235, 14)    <= sub_wire22(14);
	sub_wire2(235, 15)    <= sub_wire22(15);
	sub_wire2(235, 16)    <= sub_wire22(16);
	sub_wire2(235, 17)    <= sub_wire22(17);
	sub_wire2(235, 18)    <= sub_wire22(18);
	sub_wire2(235, 19)    <= sub_wire22(19);
	sub_wire2(235, 20)    <= sub_wire22(20);
	sub_wire2(235, 21)    <= sub_wire22(21);
	sub_wire2(235, 22)    <= sub_wire22(22);
	sub_wire2(235, 23)    <= sub_wire22(23);
	sub_wire2(235, 24)    <= sub_wire22(24);
	sub_wire2(235, 25)    <= sub_wire22(25);
	sub_wire2(235, 26)    <= sub_wire22(26);
	sub_wire2(235, 27)    <= sub_wire22(27);
	sub_wire2(235, 28)    <= sub_wire22(28);
	sub_wire2(235, 29)    <= sub_wire22(29);
	sub_wire2(235, 30)    <= sub_wire22(30);
	sub_wire2(235, 31)    <= sub_wire22(31);
	sub_wire2(235, 32)    <= sub_wire22(32);
	sub_wire2(235, 33)    <= sub_wire22(33);
	sub_wire2(235, 34)    <= sub_wire22(34);
	sub_wire2(235, 35)    <= sub_wire22(35);
	sub_wire2(235, 36)    <= sub_wire22(36);
	sub_wire2(235, 37)    <= sub_wire22(37);
	sub_wire2(235, 38)    <= sub_wire22(38);
	sub_wire2(235, 39)    <= sub_wire22(39);
	sub_wire2(234, 0)    <= sub_wire23(0);
	sub_wire2(234, 1)    <= sub_wire23(1);
	sub_wire2(234, 2)    <= sub_wire23(2);
	sub_wire2(234, 3)    <= sub_wire23(3);
	sub_wire2(234, 4)    <= sub_wire23(4);
	sub_wire2(234, 5)    <= sub_wire23(5);
	sub_wire2(234, 6)    <= sub_wire23(6);
	sub_wire2(234, 7)    <= sub_wire23(7);
	sub_wire2(234, 8)    <= sub_wire23(8);
	sub_wire2(234, 9)    <= sub_wire23(9);
	sub_wire2(234, 10)    <= sub_wire23(10);
	sub_wire2(234, 11)    <= sub_wire23(11);
	sub_wire2(234, 12)    <= sub_wire23(12);
	sub_wire2(234, 13)    <= sub_wire23(13);
	sub_wire2(234, 14)    <= sub_wire23(14);
	sub_wire2(234, 15)    <= sub_wire23(15);
	sub_wire2(234, 16)    <= sub_wire23(16);
	sub_wire2(234, 17)    <= sub_wire23(17);
	sub_wire2(234, 18)    <= sub_wire23(18);
	sub_wire2(234, 19)    <= sub_wire23(19);
	sub_wire2(234, 20)    <= sub_wire23(20);
	sub_wire2(234, 21)    <= sub_wire23(21);
	sub_wire2(234, 22)    <= sub_wire23(22);
	sub_wire2(234, 23)    <= sub_wire23(23);
	sub_wire2(234, 24)    <= sub_wire23(24);
	sub_wire2(234, 25)    <= sub_wire23(25);
	sub_wire2(234, 26)    <= sub_wire23(26);
	sub_wire2(234, 27)    <= sub_wire23(27);
	sub_wire2(234, 28)    <= sub_wire23(28);
	sub_wire2(234, 29)    <= sub_wire23(29);
	sub_wire2(234, 30)    <= sub_wire23(30);
	sub_wire2(234, 31)    <= sub_wire23(31);
	sub_wire2(234, 32)    <= sub_wire23(32);
	sub_wire2(234, 33)    <= sub_wire23(33);
	sub_wire2(234, 34)    <= sub_wire23(34);
	sub_wire2(234, 35)    <= sub_wire23(35);
	sub_wire2(234, 36)    <= sub_wire23(36);
	sub_wire2(234, 37)    <= sub_wire23(37);
	sub_wire2(234, 38)    <= sub_wire23(38);
	sub_wire2(234, 39)    <= sub_wire23(39);
	sub_wire2(233, 0)    <= sub_wire24(0);
	sub_wire2(233, 1)    <= sub_wire24(1);
	sub_wire2(233, 2)    <= sub_wire24(2);
	sub_wire2(233, 3)    <= sub_wire24(3);
	sub_wire2(233, 4)    <= sub_wire24(4);
	sub_wire2(233, 5)    <= sub_wire24(5);
	sub_wire2(233, 6)    <= sub_wire24(6);
	sub_wire2(233, 7)    <= sub_wire24(7);
	sub_wire2(233, 8)    <= sub_wire24(8);
	sub_wire2(233, 9)    <= sub_wire24(9);
	sub_wire2(233, 10)    <= sub_wire24(10);
	sub_wire2(233, 11)    <= sub_wire24(11);
	sub_wire2(233, 12)    <= sub_wire24(12);
	sub_wire2(233, 13)    <= sub_wire24(13);
	sub_wire2(233, 14)    <= sub_wire24(14);
	sub_wire2(233, 15)    <= sub_wire24(15);
	sub_wire2(233, 16)    <= sub_wire24(16);
	sub_wire2(233, 17)    <= sub_wire24(17);
	sub_wire2(233, 18)    <= sub_wire24(18);
	sub_wire2(233, 19)    <= sub_wire24(19);
	sub_wire2(233, 20)    <= sub_wire24(20);
	sub_wire2(233, 21)    <= sub_wire24(21);
	sub_wire2(233, 22)    <= sub_wire24(22);
	sub_wire2(233, 23)    <= sub_wire24(23);
	sub_wire2(233, 24)    <= sub_wire24(24);
	sub_wire2(233, 25)    <= sub_wire24(25);
	sub_wire2(233, 26)    <= sub_wire24(26);
	sub_wire2(233, 27)    <= sub_wire24(27);
	sub_wire2(233, 28)    <= sub_wire24(28);
	sub_wire2(233, 29)    <= sub_wire24(29);
	sub_wire2(233, 30)    <= sub_wire24(30);
	sub_wire2(233, 31)    <= sub_wire24(31);
	sub_wire2(233, 32)    <= sub_wire24(32);
	sub_wire2(233, 33)    <= sub_wire24(33);
	sub_wire2(233, 34)    <= sub_wire24(34);
	sub_wire2(233, 35)    <= sub_wire24(35);
	sub_wire2(233, 36)    <= sub_wire24(36);
	sub_wire2(233, 37)    <= sub_wire24(37);
	sub_wire2(233, 38)    <= sub_wire24(38);
	sub_wire2(233, 39)    <= sub_wire24(39);
	sub_wire2(232, 0)    <= sub_wire25(0);
	sub_wire2(232, 1)    <= sub_wire25(1);
	sub_wire2(232, 2)    <= sub_wire25(2);
	sub_wire2(232, 3)    <= sub_wire25(3);
	sub_wire2(232, 4)    <= sub_wire25(4);
	sub_wire2(232, 5)    <= sub_wire25(5);
	sub_wire2(232, 6)    <= sub_wire25(6);
	sub_wire2(232, 7)    <= sub_wire25(7);
	sub_wire2(232, 8)    <= sub_wire25(8);
	sub_wire2(232, 9)    <= sub_wire25(9);
	sub_wire2(232, 10)    <= sub_wire25(10);
	sub_wire2(232, 11)    <= sub_wire25(11);
	sub_wire2(232, 12)    <= sub_wire25(12);
	sub_wire2(232, 13)    <= sub_wire25(13);
	sub_wire2(232, 14)    <= sub_wire25(14);
	sub_wire2(232, 15)    <= sub_wire25(15);
	sub_wire2(232, 16)    <= sub_wire25(16);
	sub_wire2(232, 17)    <= sub_wire25(17);
	sub_wire2(232, 18)    <= sub_wire25(18);
	sub_wire2(232, 19)    <= sub_wire25(19);
	sub_wire2(232, 20)    <= sub_wire25(20);
	sub_wire2(232, 21)    <= sub_wire25(21);
	sub_wire2(232, 22)    <= sub_wire25(22);
	sub_wire2(232, 23)    <= sub_wire25(23);
	sub_wire2(232, 24)    <= sub_wire25(24);
	sub_wire2(232, 25)    <= sub_wire25(25);
	sub_wire2(232, 26)    <= sub_wire25(26);
	sub_wire2(232, 27)    <= sub_wire25(27);
	sub_wire2(232, 28)    <= sub_wire25(28);
	sub_wire2(232, 29)    <= sub_wire25(29);
	sub_wire2(232, 30)    <= sub_wire25(30);
	sub_wire2(232, 31)    <= sub_wire25(31);
	sub_wire2(232, 32)    <= sub_wire25(32);
	sub_wire2(232, 33)    <= sub_wire25(33);
	sub_wire2(232, 34)    <= sub_wire25(34);
	sub_wire2(232, 35)    <= sub_wire25(35);
	sub_wire2(232, 36)    <= sub_wire25(36);
	sub_wire2(232, 37)    <= sub_wire25(37);
	sub_wire2(232, 38)    <= sub_wire25(38);
	sub_wire2(232, 39)    <= sub_wire25(39);
	sub_wire2(231, 0)    <= sub_wire26(0);
	sub_wire2(231, 1)    <= sub_wire26(1);
	sub_wire2(231, 2)    <= sub_wire26(2);
	sub_wire2(231, 3)    <= sub_wire26(3);
	sub_wire2(231, 4)    <= sub_wire26(4);
	sub_wire2(231, 5)    <= sub_wire26(5);
	sub_wire2(231, 6)    <= sub_wire26(6);
	sub_wire2(231, 7)    <= sub_wire26(7);
	sub_wire2(231, 8)    <= sub_wire26(8);
	sub_wire2(231, 9)    <= sub_wire26(9);
	sub_wire2(231, 10)    <= sub_wire26(10);
	sub_wire2(231, 11)    <= sub_wire26(11);
	sub_wire2(231, 12)    <= sub_wire26(12);
	sub_wire2(231, 13)    <= sub_wire26(13);
	sub_wire2(231, 14)    <= sub_wire26(14);
	sub_wire2(231, 15)    <= sub_wire26(15);
	sub_wire2(231, 16)    <= sub_wire26(16);
	sub_wire2(231, 17)    <= sub_wire26(17);
	sub_wire2(231, 18)    <= sub_wire26(18);
	sub_wire2(231, 19)    <= sub_wire26(19);
	sub_wire2(231, 20)    <= sub_wire26(20);
	sub_wire2(231, 21)    <= sub_wire26(21);
	sub_wire2(231, 22)    <= sub_wire26(22);
	sub_wire2(231, 23)    <= sub_wire26(23);
	sub_wire2(231, 24)    <= sub_wire26(24);
	sub_wire2(231, 25)    <= sub_wire26(25);
	sub_wire2(231, 26)    <= sub_wire26(26);
	sub_wire2(231, 27)    <= sub_wire26(27);
	sub_wire2(231, 28)    <= sub_wire26(28);
	sub_wire2(231, 29)    <= sub_wire26(29);
	sub_wire2(231, 30)    <= sub_wire26(30);
	sub_wire2(231, 31)    <= sub_wire26(31);
	sub_wire2(231, 32)    <= sub_wire26(32);
	sub_wire2(231, 33)    <= sub_wire26(33);
	sub_wire2(231, 34)    <= sub_wire26(34);
	sub_wire2(231, 35)    <= sub_wire26(35);
	sub_wire2(231, 36)    <= sub_wire26(36);
	sub_wire2(231, 37)    <= sub_wire26(37);
	sub_wire2(231, 38)    <= sub_wire26(38);
	sub_wire2(231, 39)    <= sub_wire26(39);
	sub_wire2(230, 0)    <= sub_wire27(0);
	sub_wire2(230, 1)    <= sub_wire27(1);
	sub_wire2(230, 2)    <= sub_wire27(2);
	sub_wire2(230, 3)    <= sub_wire27(3);
	sub_wire2(230, 4)    <= sub_wire27(4);
	sub_wire2(230, 5)    <= sub_wire27(5);
	sub_wire2(230, 6)    <= sub_wire27(6);
	sub_wire2(230, 7)    <= sub_wire27(7);
	sub_wire2(230, 8)    <= sub_wire27(8);
	sub_wire2(230, 9)    <= sub_wire27(9);
	sub_wire2(230, 10)    <= sub_wire27(10);
	sub_wire2(230, 11)    <= sub_wire27(11);
	sub_wire2(230, 12)    <= sub_wire27(12);
	sub_wire2(230, 13)    <= sub_wire27(13);
	sub_wire2(230, 14)    <= sub_wire27(14);
	sub_wire2(230, 15)    <= sub_wire27(15);
	sub_wire2(230, 16)    <= sub_wire27(16);
	sub_wire2(230, 17)    <= sub_wire27(17);
	sub_wire2(230, 18)    <= sub_wire27(18);
	sub_wire2(230, 19)    <= sub_wire27(19);
	sub_wire2(230, 20)    <= sub_wire27(20);
	sub_wire2(230, 21)    <= sub_wire27(21);
	sub_wire2(230, 22)    <= sub_wire27(22);
	sub_wire2(230, 23)    <= sub_wire27(23);
	sub_wire2(230, 24)    <= sub_wire27(24);
	sub_wire2(230, 25)    <= sub_wire27(25);
	sub_wire2(230, 26)    <= sub_wire27(26);
	sub_wire2(230, 27)    <= sub_wire27(27);
	sub_wire2(230, 28)    <= sub_wire27(28);
	sub_wire2(230, 29)    <= sub_wire27(29);
	sub_wire2(230, 30)    <= sub_wire27(30);
	sub_wire2(230, 31)    <= sub_wire27(31);
	sub_wire2(230, 32)    <= sub_wire27(32);
	sub_wire2(230, 33)    <= sub_wire27(33);
	sub_wire2(230, 34)    <= sub_wire27(34);
	sub_wire2(230, 35)    <= sub_wire27(35);
	sub_wire2(230, 36)    <= sub_wire27(36);
	sub_wire2(230, 37)    <= sub_wire27(37);
	sub_wire2(230, 38)    <= sub_wire27(38);
	sub_wire2(230, 39)    <= sub_wire27(39);
	sub_wire2(229, 0)    <= sub_wire28(0);
	sub_wire2(229, 1)    <= sub_wire28(1);
	sub_wire2(229, 2)    <= sub_wire28(2);
	sub_wire2(229, 3)    <= sub_wire28(3);
	sub_wire2(229, 4)    <= sub_wire28(4);
	sub_wire2(229, 5)    <= sub_wire28(5);
	sub_wire2(229, 6)    <= sub_wire28(6);
	sub_wire2(229, 7)    <= sub_wire28(7);
	sub_wire2(229, 8)    <= sub_wire28(8);
	sub_wire2(229, 9)    <= sub_wire28(9);
	sub_wire2(229, 10)    <= sub_wire28(10);
	sub_wire2(229, 11)    <= sub_wire28(11);
	sub_wire2(229, 12)    <= sub_wire28(12);
	sub_wire2(229, 13)    <= sub_wire28(13);
	sub_wire2(229, 14)    <= sub_wire28(14);
	sub_wire2(229, 15)    <= sub_wire28(15);
	sub_wire2(229, 16)    <= sub_wire28(16);
	sub_wire2(229, 17)    <= sub_wire28(17);
	sub_wire2(229, 18)    <= sub_wire28(18);
	sub_wire2(229, 19)    <= sub_wire28(19);
	sub_wire2(229, 20)    <= sub_wire28(20);
	sub_wire2(229, 21)    <= sub_wire28(21);
	sub_wire2(229, 22)    <= sub_wire28(22);
	sub_wire2(229, 23)    <= sub_wire28(23);
	sub_wire2(229, 24)    <= sub_wire28(24);
	sub_wire2(229, 25)    <= sub_wire28(25);
	sub_wire2(229, 26)    <= sub_wire28(26);
	sub_wire2(229, 27)    <= sub_wire28(27);
	sub_wire2(229, 28)    <= sub_wire28(28);
	sub_wire2(229, 29)    <= sub_wire28(29);
	sub_wire2(229, 30)    <= sub_wire28(30);
	sub_wire2(229, 31)    <= sub_wire28(31);
	sub_wire2(229, 32)    <= sub_wire28(32);
	sub_wire2(229, 33)    <= sub_wire28(33);
	sub_wire2(229, 34)    <= sub_wire28(34);
	sub_wire2(229, 35)    <= sub_wire28(35);
	sub_wire2(229, 36)    <= sub_wire28(36);
	sub_wire2(229, 37)    <= sub_wire28(37);
	sub_wire2(229, 38)    <= sub_wire28(38);
	sub_wire2(229, 39)    <= sub_wire28(39);
	sub_wire2(228, 0)    <= sub_wire29(0);
	sub_wire2(228, 1)    <= sub_wire29(1);
	sub_wire2(228, 2)    <= sub_wire29(2);
	sub_wire2(228, 3)    <= sub_wire29(3);
	sub_wire2(228, 4)    <= sub_wire29(4);
	sub_wire2(228, 5)    <= sub_wire29(5);
	sub_wire2(228, 6)    <= sub_wire29(6);
	sub_wire2(228, 7)    <= sub_wire29(7);
	sub_wire2(228, 8)    <= sub_wire29(8);
	sub_wire2(228, 9)    <= sub_wire29(9);
	sub_wire2(228, 10)    <= sub_wire29(10);
	sub_wire2(228, 11)    <= sub_wire29(11);
	sub_wire2(228, 12)    <= sub_wire29(12);
	sub_wire2(228, 13)    <= sub_wire29(13);
	sub_wire2(228, 14)    <= sub_wire29(14);
	sub_wire2(228, 15)    <= sub_wire29(15);
	sub_wire2(228, 16)    <= sub_wire29(16);
	sub_wire2(228, 17)    <= sub_wire29(17);
	sub_wire2(228, 18)    <= sub_wire29(18);
	sub_wire2(228, 19)    <= sub_wire29(19);
	sub_wire2(228, 20)    <= sub_wire29(20);
	sub_wire2(228, 21)    <= sub_wire29(21);
	sub_wire2(228, 22)    <= sub_wire29(22);
	sub_wire2(228, 23)    <= sub_wire29(23);
	sub_wire2(228, 24)    <= sub_wire29(24);
	sub_wire2(228, 25)    <= sub_wire29(25);
	sub_wire2(228, 26)    <= sub_wire29(26);
	sub_wire2(228, 27)    <= sub_wire29(27);
	sub_wire2(228, 28)    <= sub_wire29(28);
	sub_wire2(228, 29)    <= sub_wire29(29);
	sub_wire2(228, 30)    <= sub_wire29(30);
	sub_wire2(228, 31)    <= sub_wire29(31);
	sub_wire2(228, 32)    <= sub_wire29(32);
	sub_wire2(228, 33)    <= sub_wire29(33);
	sub_wire2(228, 34)    <= sub_wire29(34);
	sub_wire2(228, 35)    <= sub_wire29(35);
	sub_wire2(228, 36)    <= sub_wire29(36);
	sub_wire2(228, 37)    <= sub_wire29(37);
	sub_wire2(228, 38)    <= sub_wire29(38);
	sub_wire2(228, 39)    <= sub_wire29(39);
	sub_wire2(227, 0)    <= sub_wire30(0);
	sub_wire2(227, 1)    <= sub_wire30(1);
	sub_wire2(227, 2)    <= sub_wire30(2);
	sub_wire2(227, 3)    <= sub_wire30(3);
	sub_wire2(227, 4)    <= sub_wire30(4);
	sub_wire2(227, 5)    <= sub_wire30(5);
	sub_wire2(227, 6)    <= sub_wire30(6);
	sub_wire2(227, 7)    <= sub_wire30(7);
	sub_wire2(227, 8)    <= sub_wire30(8);
	sub_wire2(227, 9)    <= sub_wire30(9);
	sub_wire2(227, 10)    <= sub_wire30(10);
	sub_wire2(227, 11)    <= sub_wire30(11);
	sub_wire2(227, 12)    <= sub_wire30(12);
	sub_wire2(227, 13)    <= sub_wire30(13);
	sub_wire2(227, 14)    <= sub_wire30(14);
	sub_wire2(227, 15)    <= sub_wire30(15);
	sub_wire2(227, 16)    <= sub_wire30(16);
	sub_wire2(227, 17)    <= sub_wire30(17);
	sub_wire2(227, 18)    <= sub_wire30(18);
	sub_wire2(227, 19)    <= sub_wire30(19);
	sub_wire2(227, 20)    <= sub_wire30(20);
	sub_wire2(227, 21)    <= sub_wire30(21);
	sub_wire2(227, 22)    <= sub_wire30(22);
	sub_wire2(227, 23)    <= sub_wire30(23);
	sub_wire2(227, 24)    <= sub_wire30(24);
	sub_wire2(227, 25)    <= sub_wire30(25);
	sub_wire2(227, 26)    <= sub_wire30(26);
	sub_wire2(227, 27)    <= sub_wire30(27);
	sub_wire2(227, 28)    <= sub_wire30(28);
	sub_wire2(227, 29)    <= sub_wire30(29);
	sub_wire2(227, 30)    <= sub_wire30(30);
	sub_wire2(227, 31)    <= sub_wire30(31);
	sub_wire2(227, 32)    <= sub_wire30(32);
	sub_wire2(227, 33)    <= sub_wire30(33);
	sub_wire2(227, 34)    <= sub_wire30(34);
	sub_wire2(227, 35)    <= sub_wire30(35);
	sub_wire2(227, 36)    <= sub_wire30(36);
	sub_wire2(227, 37)    <= sub_wire30(37);
	sub_wire2(227, 38)    <= sub_wire30(38);
	sub_wire2(227, 39)    <= sub_wire30(39);
	sub_wire2(226, 0)    <= sub_wire31(0);
	sub_wire2(226, 1)    <= sub_wire31(1);
	sub_wire2(226, 2)    <= sub_wire31(2);
	sub_wire2(226, 3)    <= sub_wire31(3);
	sub_wire2(226, 4)    <= sub_wire31(4);
	sub_wire2(226, 5)    <= sub_wire31(5);
	sub_wire2(226, 6)    <= sub_wire31(6);
	sub_wire2(226, 7)    <= sub_wire31(7);
	sub_wire2(226, 8)    <= sub_wire31(8);
	sub_wire2(226, 9)    <= sub_wire31(9);
	sub_wire2(226, 10)    <= sub_wire31(10);
	sub_wire2(226, 11)    <= sub_wire31(11);
	sub_wire2(226, 12)    <= sub_wire31(12);
	sub_wire2(226, 13)    <= sub_wire31(13);
	sub_wire2(226, 14)    <= sub_wire31(14);
	sub_wire2(226, 15)    <= sub_wire31(15);
	sub_wire2(226, 16)    <= sub_wire31(16);
	sub_wire2(226, 17)    <= sub_wire31(17);
	sub_wire2(226, 18)    <= sub_wire31(18);
	sub_wire2(226, 19)    <= sub_wire31(19);
	sub_wire2(226, 20)    <= sub_wire31(20);
	sub_wire2(226, 21)    <= sub_wire31(21);
	sub_wire2(226, 22)    <= sub_wire31(22);
	sub_wire2(226, 23)    <= sub_wire31(23);
	sub_wire2(226, 24)    <= sub_wire31(24);
	sub_wire2(226, 25)    <= sub_wire31(25);
	sub_wire2(226, 26)    <= sub_wire31(26);
	sub_wire2(226, 27)    <= sub_wire31(27);
	sub_wire2(226, 28)    <= sub_wire31(28);
	sub_wire2(226, 29)    <= sub_wire31(29);
	sub_wire2(226, 30)    <= sub_wire31(30);
	sub_wire2(226, 31)    <= sub_wire31(31);
	sub_wire2(226, 32)    <= sub_wire31(32);
	sub_wire2(226, 33)    <= sub_wire31(33);
	sub_wire2(226, 34)    <= sub_wire31(34);
	sub_wire2(226, 35)    <= sub_wire31(35);
	sub_wire2(226, 36)    <= sub_wire31(36);
	sub_wire2(226, 37)    <= sub_wire31(37);
	sub_wire2(226, 38)    <= sub_wire31(38);
	sub_wire2(226, 39)    <= sub_wire31(39);
	sub_wire2(225, 0)    <= sub_wire32(0);
	sub_wire2(225, 1)    <= sub_wire32(1);
	sub_wire2(225, 2)    <= sub_wire32(2);
	sub_wire2(225, 3)    <= sub_wire32(3);
	sub_wire2(225, 4)    <= sub_wire32(4);
	sub_wire2(225, 5)    <= sub_wire32(5);
	sub_wire2(225, 6)    <= sub_wire32(6);
	sub_wire2(225, 7)    <= sub_wire32(7);
	sub_wire2(225, 8)    <= sub_wire32(8);
	sub_wire2(225, 9)    <= sub_wire32(9);
	sub_wire2(225, 10)    <= sub_wire32(10);
	sub_wire2(225, 11)    <= sub_wire32(11);
	sub_wire2(225, 12)    <= sub_wire32(12);
	sub_wire2(225, 13)    <= sub_wire32(13);
	sub_wire2(225, 14)    <= sub_wire32(14);
	sub_wire2(225, 15)    <= sub_wire32(15);
	sub_wire2(225, 16)    <= sub_wire32(16);
	sub_wire2(225, 17)    <= sub_wire32(17);
	sub_wire2(225, 18)    <= sub_wire32(18);
	sub_wire2(225, 19)    <= sub_wire32(19);
	sub_wire2(225, 20)    <= sub_wire32(20);
	sub_wire2(225, 21)    <= sub_wire32(21);
	sub_wire2(225, 22)    <= sub_wire32(22);
	sub_wire2(225, 23)    <= sub_wire32(23);
	sub_wire2(225, 24)    <= sub_wire32(24);
	sub_wire2(225, 25)    <= sub_wire32(25);
	sub_wire2(225, 26)    <= sub_wire32(26);
	sub_wire2(225, 27)    <= sub_wire32(27);
	sub_wire2(225, 28)    <= sub_wire32(28);
	sub_wire2(225, 29)    <= sub_wire32(29);
	sub_wire2(225, 30)    <= sub_wire32(30);
	sub_wire2(225, 31)    <= sub_wire32(31);
	sub_wire2(225, 32)    <= sub_wire32(32);
	sub_wire2(225, 33)    <= sub_wire32(33);
	sub_wire2(225, 34)    <= sub_wire32(34);
	sub_wire2(225, 35)    <= sub_wire32(35);
	sub_wire2(225, 36)    <= sub_wire32(36);
	sub_wire2(225, 37)    <= sub_wire32(37);
	sub_wire2(225, 38)    <= sub_wire32(38);
	sub_wire2(225, 39)    <= sub_wire32(39);
	sub_wire2(224, 0)    <= sub_wire33(0);
	sub_wire2(224, 1)    <= sub_wire33(1);
	sub_wire2(224, 2)    <= sub_wire33(2);
	sub_wire2(224, 3)    <= sub_wire33(3);
	sub_wire2(224, 4)    <= sub_wire33(4);
	sub_wire2(224, 5)    <= sub_wire33(5);
	sub_wire2(224, 6)    <= sub_wire33(6);
	sub_wire2(224, 7)    <= sub_wire33(7);
	sub_wire2(224, 8)    <= sub_wire33(8);
	sub_wire2(224, 9)    <= sub_wire33(9);
	sub_wire2(224, 10)    <= sub_wire33(10);
	sub_wire2(224, 11)    <= sub_wire33(11);
	sub_wire2(224, 12)    <= sub_wire33(12);
	sub_wire2(224, 13)    <= sub_wire33(13);
	sub_wire2(224, 14)    <= sub_wire33(14);
	sub_wire2(224, 15)    <= sub_wire33(15);
	sub_wire2(224, 16)    <= sub_wire33(16);
	sub_wire2(224, 17)    <= sub_wire33(17);
	sub_wire2(224, 18)    <= sub_wire33(18);
	sub_wire2(224, 19)    <= sub_wire33(19);
	sub_wire2(224, 20)    <= sub_wire33(20);
	sub_wire2(224, 21)    <= sub_wire33(21);
	sub_wire2(224, 22)    <= sub_wire33(22);
	sub_wire2(224, 23)    <= sub_wire33(23);
	sub_wire2(224, 24)    <= sub_wire33(24);
	sub_wire2(224, 25)    <= sub_wire33(25);
	sub_wire2(224, 26)    <= sub_wire33(26);
	sub_wire2(224, 27)    <= sub_wire33(27);
	sub_wire2(224, 28)    <= sub_wire33(28);
	sub_wire2(224, 29)    <= sub_wire33(29);
	sub_wire2(224, 30)    <= sub_wire33(30);
	sub_wire2(224, 31)    <= sub_wire33(31);
	sub_wire2(224, 32)    <= sub_wire33(32);
	sub_wire2(224, 33)    <= sub_wire33(33);
	sub_wire2(224, 34)    <= sub_wire33(34);
	sub_wire2(224, 35)    <= sub_wire33(35);
	sub_wire2(224, 36)    <= sub_wire33(36);
	sub_wire2(224, 37)    <= sub_wire33(37);
	sub_wire2(224, 38)    <= sub_wire33(38);
	sub_wire2(224, 39)    <= sub_wire33(39);
	sub_wire2(223, 0)    <= sub_wire34(0);
	sub_wire2(223, 1)    <= sub_wire34(1);
	sub_wire2(223, 2)    <= sub_wire34(2);
	sub_wire2(223, 3)    <= sub_wire34(3);
	sub_wire2(223, 4)    <= sub_wire34(4);
	sub_wire2(223, 5)    <= sub_wire34(5);
	sub_wire2(223, 6)    <= sub_wire34(6);
	sub_wire2(223, 7)    <= sub_wire34(7);
	sub_wire2(223, 8)    <= sub_wire34(8);
	sub_wire2(223, 9)    <= sub_wire34(9);
	sub_wire2(223, 10)    <= sub_wire34(10);
	sub_wire2(223, 11)    <= sub_wire34(11);
	sub_wire2(223, 12)    <= sub_wire34(12);
	sub_wire2(223, 13)    <= sub_wire34(13);
	sub_wire2(223, 14)    <= sub_wire34(14);
	sub_wire2(223, 15)    <= sub_wire34(15);
	sub_wire2(223, 16)    <= sub_wire34(16);
	sub_wire2(223, 17)    <= sub_wire34(17);
	sub_wire2(223, 18)    <= sub_wire34(18);
	sub_wire2(223, 19)    <= sub_wire34(19);
	sub_wire2(223, 20)    <= sub_wire34(20);
	sub_wire2(223, 21)    <= sub_wire34(21);
	sub_wire2(223, 22)    <= sub_wire34(22);
	sub_wire2(223, 23)    <= sub_wire34(23);
	sub_wire2(223, 24)    <= sub_wire34(24);
	sub_wire2(223, 25)    <= sub_wire34(25);
	sub_wire2(223, 26)    <= sub_wire34(26);
	sub_wire2(223, 27)    <= sub_wire34(27);
	sub_wire2(223, 28)    <= sub_wire34(28);
	sub_wire2(223, 29)    <= sub_wire34(29);
	sub_wire2(223, 30)    <= sub_wire34(30);
	sub_wire2(223, 31)    <= sub_wire34(31);
	sub_wire2(223, 32)    <= sub_wire34(32);
	sub_wire2(223, 33)    <= sub_wire34(33);
	sub_wire2(223, 34)    <= sub_wire34(34);
	sub_wire2(223, 35)    <= sub_wire34(35);
	sub_wire2(223, 36)    <= sub_wire34(36);
	sub_wire2(223, 37)    <= sub_wire34(37);
	sub_wire2(223, 38)    <= sub_wire34(38);
	sub_wire2(223, 39)    <= sub_wire34(39);
	sub_wire2(222, 0)    <= sub_wire35(0);
	sub_wire2(222, 1)    <= sub_wire35(1);
	sub_wire2(222, 2)    <= sub_wire35(2);
	sub_wire2(222, 3)    <= sub_wire35(3);
	sub_wire2(222, 4)    <= sub_wire35(4);
	sub_wire2(222, 5)    <= sub_wire35(5);
	sub_wire2(222, 6)    <= sub_wire35(6);
	sub_wire2(222, 7)    <= sub_wire35(7);
	sub_wire2(222, 8)    <= sub_wire35(8);
	sub_wire2(222, 9)    <= sub_wire35(9);
	sub_wire2(222, 10)    <= sub_wire35(10);
	sub_wire2(222, 11)    <= sub_wire35(11);
	sub_wire2(222, 12)    <= sub_wire35(12);
	sub_wire2(222, 13)    <= sub_wire35(13);
	sub_wire2(222, 14)    <= sub_wire35(14);
	sub_wire2(222, 15)    <= sub_wire35(15);
	sub_wire2(222, 16)    <= sub_wire35(16);
	sub_wire2(222, 17)    <= sub_wire35(17);
	sub_wire2(222, 18)    <= sub_wire35(18);
	sub_wire2(222, 19)    <= sub_wire35(19);
	sub_wire2(222, 20)    <= sub_wire35(20);
	sub_wire2(222, 21)    <= sub_wire35(21);
	sub_wire2(222, 22)    <= sub_wire35(22);
	sub_wire2(222, 23)    <= sub_wire35(23);
	sub_wire2(222, 24)    <= sub_wire35(24);
	sub_wire2(222, 25)    <= sub_wire35(25);
	sub_wire2(222, 26)    <= sub_wire35(26);
	sub_wire2(222, 27)    <= sub_wire35(27);
	sub_wire2(222, 28)    <= sub_wire35(28);
	sub_wire2(222, 29)    <= sub_wire35(29);
	sub_wire2(222, 30)    <= sub_wire35(30);
	sub_wire2(222, 31)    <= sub_wire35(31);
	sub_wire2(222, 32)    <= sub_wire35(32);
	sub_wire2(222, 33)    <= sub_wire35(33);
	sub_wire2(222, 34)    <= sub_wire35(34);
	sub_wire2(222, 35)    <= sub_wire35(35);
	sub_wire2(222, 36)    <= sub_wire35(36);
	sub_wire2(222, 37)    <= sub_wire35(37);
	sub_wire2(222, 38)    <= sub_wire35(38);
	sub_wire2(222, 39)    <= sub_wire35(39);
	sub_wire2(221, 0)    <= sub_wire36(0);
	sub_wire2(221, 1)    <= sub_wire36(1);
	sub_wire2(221, 2)    <= sub_wire36(2);
	sub_wire2(221, 3)    <= sub_wire36(3);
	sub_wire2(221, 4)    <= sub_wire36(4);
	sub_wire2(221, 5)    <= sub_wire36(5);
	sub_wire2(221, 6)    <= sub_wire36(6);
	sub_wire2(221, 7)    <= sub_wire36(7);
	sub_wire2(221, 8)    <= sub_wire36(8);
	sub_wire2(221, 9)    <= sub_wire36(9);
	sub_wire2(221, 10)    <= sub_wire36(10);
	sub_wire2(221, 11)    <= sub_wire36(11);
	sub_wire2(221, 12)    <= sub_wire36(12);
	sub_wire2(221, 13)    <= sub_wire36(13);
	sub_wire2(221, 14)    <= sub_wire36(14);
	sub_wire2(221, 15)    <= sub_wire36(15);
	sub_wire2(221, 16)    <= sub_wire36(16);
	sub_wire2(221, 17)    <= sub_wire36(17);
	sub_wire2(221, 18)    <= sub_wire36(18);
	sub_wire2(221, 19)    <= sub_wire36(19);
	sub_wire2(221, 20)    <= sub_wire36(20);
	sub_wire2(221, 21)    <= sub_wire36(21);
	sub_wire2(221, 22)    <= sub_wire36(22);
	sub_wire2(221, 23)    <= sub_wire36(23);
	sub_wire2(221, 24)    <= sub_wire36(24);
	sub_wire2(221, 25)    <= sub_wire36(25);
	sub_wire2(221, 26)    <= sub_wire36(26);
	sub_wire2(221, 27)    <= sub_wire36(27);
	sub_wire2(221, 28)    <= sub_wire36(28);
	sub_wire2(221, 29)    <= sub_wire36(29);
	sub_wire2(221, 30)    <= sub_wire36(30);
	sub_wire2(221, 31)    <= sub_wire36(31);
	sub_wire2(221, 32)    <= sub_wire36(32);
	sub_wire2(221, 33)    <= sub_wire36(33);
	sub_wire2(221, 34)    <= sub_wire36(34);
	sub_wire2(221, 35)    <= sub_wire36(35);
	sub_wire2(221, 36)    <= sub_wire36(36);
	sub_wire2(221, 37)    <= sub_wire36(37);
	sub_wire2(221, 38)    <= sub_wire36(38);
	sub_wire2(221, 39)    <= sub_wire36(39);
	sub_wire2(220, 0)    <= sub_wire37(0);
	sub_wire2(220, 1)    <= sub_wire37(1);
	sub_wire2(220, 2)    <= sub_wire37(2);
	sub_wire2(220, 3)    <= sub_wire37(3);
	sub_wire2(220, 4)    <= sub_wire37(4);
	sub_wire2(220, 5)    <= sub_wire37(5);
	sub_wire2(220, 6)    <= sub_wire37(6);
	sub_wire2(220, 7)    <= sub_wire37(7);
	sub_wire2(220, 8)    <= sub_wire37(8);
	sub_wire2(220, 9)    <= sub_wire37(9);
	sub_wire2(220, 10)    <= sub_wire37(10);
	sub_wire2(220, 11)    <= sub_wire37(11);
	sub_wire2(220, 12)    <= sub_wire37(12);
	sub_wire2(220, 13)    <= sub_wire37(13);
	sub_wire2(220, 14)    <= sub_wire37(14);
	sub_wire2(220, 15)    <= sub_wire37(15);
	sub_wire2(220, 16)    <= sub_wire37(16);
	sub_wire2(220, 17)    <= sub_wire37(17);
	sub_wire2(220, 18)    <= sub_wire37(18);
	sub_wire2(220, 19)    <= sub_wire37(19);
	sub_wire2(220, 20)    <= sub_wire37(20);
	sub_wire2(220, 21)    <= sub_wire37(21);
	sub_wire2(220, 22)    <= sub_wire37(22);
	sub_wire2(220, 23)    <= sub_wire37(23);
	sub_wire2(220, 24)    <= sub_wire37(24);
	sub_wire2(220, 25)    <= sub_wire37(25);
	sub_wire2(220, 26)    <= sub_wire37(26);
	sub_wire2(220, 27)    <= sub_wire37(27);
	sub_wire2(220, 28)    <= sub_wire37(28);
	sub_wire2(220, 29)    <= sub_wire37(29);
	sub_wire2(220, 30)    <= sub_wire37(30);
	sub_wire2(220, 31)    <= sub_wire37(31);
	sub_wire2(220, 32)    <= sub_wire37(32);
	sub_wire2(220, 33)    <= sub_wire37(33);
	sub_wire2(220, 34)    <= sub_wire37(34);
	sub_wire2(220, 35)    <= sub_wire37(35);
	sub_wire2(220, 36)    <= sub_wire37(36);
	sub_wire2(220, 37)    <= sub_wire37(37);
	sub_wire2(220, 38)    <= sub_wire37(38);
	sub_wire2(220, 39)    <= sub_wire37(39);
	sub_wire2(219, 0)    <= sub_wire38(0);
	sub_wire2(219, 1)    <= sub_wire38(1);
	sub_wire2(219, 2)    <= sub_wire38(2);
	sub_wire2(219, 3)    <= sub_wire38(3);
	sub_wire2(219, 4)    <= sub_wire38(4);
	sub_wire2(219, 5)    <= sub_wire38(5);
	sub_wire2(219, 6)    <= sub_wire38(6);
	sub_wire2(219, 7)    <= sub_wire38(7);
	sub_wire2(219, 8)    <= sub_wire38(8);
	sub_wire2(219, 9)    <= sub_wire38(9);
	sub_wire2(219, 10)    <= sub_wire38(10);
	sub_wire2(219, 11)    <= sub_wire38(11);
	sub_wire2(219, 12)    <= sub_wire38(12);
	sub_wire2(219, 13)    <= sub_wire38(13);
	sub_wire2(219, 14)    <= sub_wire38(14);
	sub_wire2(219, 15)    <= sub_wire38(15);
	sub_wire2(219, 16)    <= sub_wire38(16);
	sub_wire2(219, 17)    <= sub_wire38(17);
	sub_wire2(219, 18)    <= sub_wire38(18);
	sub_wire2(219, 19)    <= sub_wire38(19);
	sub_wire2(219, 20)    <= sub_wire38(20);
	sub_wire2(219, 21)    <= sub_wire38(21);
	sub_wire2(219, 22)    <= sub_wire38(22);
	sub_wire2(219, 23)    <= sub_wire38(23);
	sub_wire2(219, 24)    <= sub_wire38(24);
	sub_wire2(219, 25)    <= sub_wire38(25);
	sub_wire2(219, 26)    <= sub_wire38(26);
	sub_wire2(219, 27)    <= sub_wire38(27);
	sub_wire2(219, 28)    <= sub_wire38(28);
	sub_wire2(219, 29)    <= sub_wire38(29);
	sub_wire2(219, 30)    <= sub_wire38(30);
	sub_wire2(219, 31)    <= sub_wire38(31);
	sub_wire2(219, 32)    <= sub_wire38(32);
	sub_wire2(219, 33)    <= sub_wire38(33);
	sub_wire2(219, 34)    <= sub_wire38(34);
	sub_wire2(219, 35)    <= sub_wire38(35);
	sub_wire2(219, 36)    <= sub_wire38(36);
	sub_wire2(219, 37)    <= sub_wire38(37);
	sub_wire2(219, 38)    <= sub_wire38(38);
	sub_wire2(219, 39)    <= sub_wire38(39);
	sub_wire2(218, 0)    <= sub_wire39(0);
	sub_wire2(218, 1)    <= sub_wire39(1);
	sub_wire2(218, 2)    <= sub_wire39(2);
	sub_wire2(218, 3)    <= sub_wire39(3);
	sub_wire2(218, 4)    <= sub_wire39(4);
	sub_wire2(218, 5)    <= sub_wire39(5);
	sub_wire2(218, 6)    <= sub_wire39(6);
	sub_wire2(218, 7)    <= sub_wire39(7);
	sub_wire2(218, 8)    <= sub_wire39(8);
	sub_wire2(218, 9)    <= sub_wire39(9);
	sub_wire2(218, 10)    <= sub_wire39(10);
	sub_wire2(218, 11)    <= sub_wire39(11);
	sub_wire2(218, 12)    <= sub_wire39(12);
	sub_wire2(218, 13)    <= sub_wire39(13);
	sub_wire2(218, 14)    <= sub_wire39(14);
	sub_wire2(218, 15)    <= sub_wire39(15);
	sub_wire2(218, 16)    <= sub_wire39(16);
	sub_wire2(218, 17)    <= sub_wire39(17);
	sub_wire2(218, 18)    <= sub_wire39(18);
	sub_wire2(218, 19)    <= sub_wire39(19);
	sub_wire2(218, 20)    <= sub_wire39(20);
	sub_wire2(218, 21)    <= sub_wire39(21);
	sub_wire2(218, 22)    <= sub_wire39(22);
	sub_wire2(218, 23)    <= sub_wire39(23);
	sub_wire2(218, 24)    <= sub_wire39(24);
	sub_wire2(218, 25)    <= sub_wire39(25);
	sub_wire2(218, 26)    <= sub_wire39(26);
	sub_wire2(218, 27)    <= sub_wire39(27);
	sub_wire2(218, 28)    <= sub_wire39(28);
	sub_wire2(218, 29)    <= sub_wire39(29);
	sub_wire2(218, 30)    <= sub_wire39(30);
	sub_wire2(218, 31)    <= sub_wire39(31);
	sub_wire2(218, 32)    <= sub_wire39(32);
	sub_wire2(218, 33)    <= sub_wire39(33);
	sub_wire2(218, 34)    <= sub_wire39(34);
	sub_wire2(218, 35)    <= sub_wire39(35);
	sub_wire2(218, 36)    <= sub_wire39(36);
	sub_wire2(218, 37)    <= sub_wire39(37);
	sub_wire2(218, 38)    <= sub_wire39(38);
	sub_wire2(218, 39)    <= sub_wire39(39);
	sub_wire2(217, 0)    <= sub_wire40(0);
	sub_wire2(217, 1)    <= sub_wire40(1);
	sub_wire2(217, 2)    <= sub_wire40(2);
	sub_wire2(217, 3)    <= sub_wire40(3);
	sub_wire2(217, 4)    <= sub_wire40(4);
	sub_wire2(217, 5)    <= sub_wire40(5);
	sub_wire2(217, 6)    <= sub_wire40(6);
	sub_wire2(217, 7)    <= sub_wire40(7);
	sub_wire2(217, 8)    <= sub_wire40(8);
	sub_wire2(217, 9)    <= sub_wire40(9);
	sub_wire2(217, 10)    <= sub_wire40(10);
	sub_wire2(217, 11)    <= sub_wire40(11);
	sub_wire2(217, 12)    <= sub_wire40(12);
	sub_wire2(217, 13)    <= sub_wire40(13);
	sub_wire2(217, 14)    <= sub_wire40(14);
	sub_wire2(217, 15)    <= sub_wire40(15);
	sub_wire2(217, 16)    <= sub_wire40(16);
	sub_wire2(217, 17)    <= sub_wire40(17);
	sub_wire2(217, 18)    <= sub_wire40(18);
	sub_wire2(217, 19)    <= sub_wire40(19);
	sub_wire2(217, 20)    <= sub_wire40(20);
	sub_wire2(217, 21)    <= sub_wire40(21);
	sub_wire2(217, 22)    <= sub_wire40(22);
	sub_wire2(217, 23)    <= sub_wire40(23);
	sub_wire2(217, 24)    <= sub_wire40(24);
	sub_wire2(217, 25)    <= sub_wire40(25);
	sub_wire2(217, 26)    <= sub_wire40(26);
	sub_wire2(217, 27)    <= sub_wire40(27);
	sub_wire2(217, 28)    <= sub_wire40(28);
	sub_wire2(217, 29)    <= sub_wire40(29);
	sub_wire2(217, 30)    <= sub_wire40(30);
	sub_wire2(217, 31)    <= sub_wire40(31);
	sub_wire2(217, 32)    <= sub_wire40(32);
	sub_wire2(217, 33)    <= sub_wire40(33);
	sub_wire2(217, 34)    <= sub_wire40(34);
	sub_wire2(217, 35)    <= sub_wire40(35);
	sub_wire2(217, 36)    <= sub_wire40(36);
	sub_wire2(217, 37)    <= sub_wire40(37);
	sub_wire2(217, 38)    <= sub_wire40(38);
	sub_wire2(217, 39)    <= sub_wire40(39);
	sub_wire2(216, 0)    <= sub_wire41(0);
	sub_wire2(216, 1)    <= sub_wire41(1);
	sub_wire2(216, 2)    <= sub_wire41(2);
	sub_wire2(216, 3)    <= sub_wire41(3);
	sub_wire2(216, 4)    <= sub_wire41(4);
	sub_wire2(216, 5)    <= sub_wire41(5);
	sub_wire2(216, 6)    <= sub_wire41(6);
	sub_wire2(216, 7)    <= sub_wire41(7);
	sub_wire2(216, 8)    <= sub_wire41(8);
	sub_wire2(216, 9)    <= sub_wire41(9);
	sub_wire2(216, 10)    <= sub_wire41(10);
	sub_wire2(216, 11)    <= sub_wire41(11);
	sub_wire2(216, 12)    <= sub_wire41(12);
	sub_wire2(216, 13)    <= sub_wire41(13);
	sub_wire2(216, 14)    <= sub_wire41(14);
	sub_wire2(216, 15)    <= sub_wire41(15);
	sub_wire2(216, 16)    <= sub_wire41(16);
	sub_wire2(216, 17)    <= sub_wire41(17);
	sub_wire2(216, 18)    <= sub_wire41(18);
	sub_wire2(216, 19)    <= sub_wire41(19);
	sub_wire2(216, 20)    <= sub_wire41(20);
	sub_wire2(216, 21)    <= sub_wire41(21);
	sub_wire2(216, 22)    <= sub_wire41(22);
	sub_wire2(216, 23)    <= sub_wire41(23);
	sub_wire2(216, 24)    <= sub_wire41(24);
	sub_wire2(216, 25)    <= sub_wire41(25);
	sub_wire2(216, 26)    <= sub_wire41(26);
	sub_wire2(216, 27)    <= sub_wire41(27);
	sub_wire2(216, 28)    <= sub_wire41(28);
	sub_wire2(216, 29)    <= sub_wire41(29);
	sub_wire2(216, 30)    <= sub_wire41(30);
	sub_wire2(216, 31)    <= sub_wire41(31);
	sub_wire2(216, 32)    <= sub_wire41(32);
	sub_wire2(216, 33)    <= sub_wire41(33);
	sub_wire2(216, 34)    <= sub_wire41(34);
	sub_wire2(216, 35)    <= sub_wire41(35);
	sub_wire2(216, 36)    <= sub_wire41(36);
	sub_wire2(216, 37)    <= sub_wire41(37);
	sub_wire2(216, 38)    <= sub_wire41(38);
	sub_wire2(216, 39)    <= sub_wire41(39);
	sub_wire2(215, 0)    <= sub_wire42(0);
	sub_wire2(215, 1)    <= sub_wire42(1);
	sub_wire2(215, 2)    <= sub_wire42(2);
	sub_wire2(215, 3)    <= sub_wire42(3);
	sub_wire2(215, 4)    <= sub_wire42(4);
	sub_wire2(215, 5)    <= sub_wire42(5);
	sub_wire2(215, 6)    <= sub_wire42(6);
	sub_wire2(215, 7)    <= sub_wire42(7);
	sub_wire2(215, 8)    <= sub_wire42(8);
	sub_wire2(215, 9)    <= sub_wire42(9);
	sub_wire2(215, 10)    <= sub_wire42(10);
	sub_wire2(215, 11)    <= sub_wire42(11);
	sub_wire2(215, 12)    <= sub_wire42(12);
	sub_wire2(215, 13)    <= sub_wire42(13);
	sub_wire2(215, 14)    <= sub_wire42(14);
	sub_wire2(215, 15)    <= sub_wire42(15);
	sub_wire2(215, 16)    <= sub_wire42(16);
	sub_wire2(215, 17)    <= sub_wire42(17);
	sub_wire2(215, 18)    <= sub_wire42(18);
	sub_wire2(215, 19)    <= sub_wire42(19);
	sub_wire2(215, 20)    <= sub_wire42(20);
	sub_wire2(215, 21)    <= sub_wire42(21);
	sub_wire2(215, 22)    <= sub_wire42(22);
	sub_wire2(215, 23)    <= sub_wire42(23);
	sub_wire2(215, 24)    <= sub_wire42(24);
	sub_wire2(215, 25)    <= sub_wire42(25);
	sub_wire2(215, 26)    <= sub_wire42(26);
	sub_wire2(215, 27)    <= sub_wire42(27);
	sub_wire2(215, 28)    <= sub_wire42(28);
	sub_wire2(215, 29)    <= sub_wire42(29);
	sub_wire2(215, 30)    <= sub_wire42(30);
	sub_wire2(215, 31)    <= sub_wire42(31);
	sub_wire2(215, 32)    <= sub_wire42(32);
	sub_wire2(215, 33)    <= sub_wire42(33);
	sub_wire2(215, 34)    <= sub_wire42(34);
	sub_wire2(215, 35)    <= sub_wire42(35);
	sub_wire2(215, 36)    <= sub_wire42(36);
	sub_wire2(215, 37)    <= sub_wire42(37);
	sub_wire2(215, 38)    <= sub_wire42(38);
	sub_wire2(215, 39)    <= sub_wire42(39);
	sub_wire2(214, 0)    <= sub_wire43(0);
	sub_wire2(214, 1)    <= sub_wire43(1);
	sub_wire2(214, 2)    <= sub_wire43(2);
	sub_wire2(214, 3)    <= sub_wire43(3);
	sub_wire2(214, 4)    <= sub_wire43(4);
	sub_wire2(214, 5)    <= sub_wire43(5);
	sub_wire2(214, 6)    <= sub_wire43(6);
	sub_wire2(214, 7)    <= sub_wire43(7);
	sub_wire2(214, 8)    <= sub_wire43(8);
	sub_wire2(214, 9)    <= sub_wire43(9);
	sub_wire2(214, 10)    <= sub_wire43(10);
	sub_wire2(214, 11)    <= sub_wire43(11);
	sub_wire2(214, 12)    <= sub_wire43(12);
	sub_wire2(214, 13)    <= sub_wire43(13);
	sub_wire2(214, 14)    <= sub_wire43(14);
	sub_wire2(214, 15)    <= sub_wire43(15);
	sub_wire2(214, 16)    <= sub_wire43(16);
	sub_wire2(214, 17)    <= sub_wire43(17);
	sub_wire2(214, 18)    <= sub_wire43(18);
	sub_wire2(214, 19)    <= sub_wire43(19);
	sub_wire2(214, 20)    <= sub_wire43(20);
	sub_wire2(214, 21)    <= sub_wire43(21);
	sub_wire2(214, 22)    <= sub_wire43(22);
	sub_wire2(214, 23)    <= sub_wire43(23);
	sub_wire2(214, 24)    <= sub_wire43(24);
	sub_wire2(214, 25)    <= sub_wire43(25);
	sub_wire2(214, 26)    <= sub_wire43(26);
	sub_wire2(214, 27)    <= sub_wire43(27);
	sub_wire2(214, 28)    <= sub_wire43(28);
	sub_wire2(214, 29)    <= sub_wire43(29);
	sub_wire2(214, 30)    <= sub_wire43(30);
	sub_wire2(214, 31)    <= sub_wire43(31);
	sub_wire2(214, 32)    <= sub_wire43(32);
	sub_wire2(214, 33)    <= sub_wire43(33);
	sub_wire2(214, 34)    <= sub_wire43(34);
	sub_wire2(214, 35)    <= sub_wire43(35);
	sub_wire2(214, 36)    <= sub_wire43(36);
	sub_wire2(214, 37)    <= sub_wire43(37);
	sub_wire2(214, 38)    <= sub_wire43(38);
	sub_wire2(214, 39)    <= sub_wire43(39);
	sub_wire2(213, 0)    <= sub_wire44(0);
	sub_wire2(213, 1)    <= sub_wire44(1);
	sub_wire2(213, 2)    <= sub_wire44(2);
	sub_wire2(213, 3)    <= sub_wire44(3);
	sub_wire2(213, 4)    <= sub_wire44(4);
	sub_wire2(213, 5)    <= sub_wire44(5);
	sub_wire2(213, 6)    <= sub_wire44(6);
	sub_wire2(213, 7)    <= sub_wire44(7);
	sub_wire2(213, 8)    <= sub_wire44(8);
	sub_wire2(213, 9)    <= sub_wire44(9);
	sub_wire2(213, 10)    <= sub_wire44(10);
	sub_wire2(213, 11)    <= sub_wire44(11);
	sub_wire2(213, 12)    <= sub_wire44(12);
	sub_wire2(213, 13)    <= sub_wire44(13);
	sub_wire2(213, 14)    <= sub_wire44(14);
	sub_wire2(213, 15)    <= sub_wire44(15);
	sub_wire2(213, 16)    <= sub_wire44(16);
	sub_wire2(213, 17)    <= sub_wire44(17);
	sub_wire2(213, 18)    <= sub_wire44(18);
	sub_wire2(213, 19)    <= sub_wire44(19);
	sub_wire2(213, 20)    <= sub_wire44(20);
	sub_wire2(213, 21)    <= sub_wire44(21);
	sub_wire2(213, 22)    <= sub_wire44(22);
	sub_wire2(213, 23)    <= sub_wire44(23);
	sub_wire2(213, 24)    <= sub_wire44(24);
	sub_wire2(213, 25)    <= sub_wire44(25);
	sub_wire2(213, 26)    <= sub_wire44(26);
	sub_wire2(213, 27)    <= sub_wire44(27);
	sub_wire2(213, 28)    <= sub_wire44(28);
	sub_wire2(213, 29)    <= sub_wire44(29);
	sub_wire2(213, 30)    <= sub_wire44(30);
	sub_wire2(213, 31)    <= sub_wire44(31);
	sub_wire2(213, 32)    <= sub_wire44(32);
	sub_wire2(213, 33)    <= sub_wire44(33);
	sub_wire2(213, 34)    <= sub_wire44(34);
	sub_wire2(213, 35)    <= sub_wire44(35);
	sub_wire2(213, 36)    <= sub_wire44(36);
	sub_wire2(213, 37)    <= sub_wire44(37);
	sub_wire2(213, 38)    <= sub_wire44(38);
	sub_wire2(213, 39)    <= sub_wire44(39);
	sub_wire2(212, 0)    <= sub_wire45(0);
	sub_wire2(212, 1)    <= sub_wire45(1);
	sub_wire2(212, 2)    <= sub_wire45(2);
	sub_wire2(212, 3)    <= sub_wire45(3);
	sub_wire2(212, 4)    <= sub_wire45(4);
	sub_wire2(212, 5)    <= sub_wire45(5);
	sub_wire2(212, 6)    <= sub_wire45(6);
	sub_wire2(212, 7)    <= sub_wire45(7);
	sub_wire2(212, 8)    <= sub_wire45(8);
	sub_wire2(212, 9)    <= sub_wire45(9);
	sub_wire2(212, 10)    <= sub_wire45(10);
	sub_wire2(212, 11)    <= sub_wire45(11);
	sub_wire2(212, 12)    <= sub_wire45(12);
	sub_wire2(212, 13)    <= sub_wire45(13);
	sub_wire2(212, 14)    <= sub_wire45(14);
	sub_wire2(212, 15)    <= sub_wire45(15);
	sub_wire2(212, 16)    <= sub_wire45(16);
	sub_wire2(212, 17)    <= sub_wire45(17);
	sub_wire2(212, 18)    <= sub_wire45(18);
	sub_wire2(212, 19)    <= sub_wire45(19);
	sub_wire2(212, 20)    <= sub_wire45(20);
	sub_wire2(212, 21)    <= sub_wire45(21);
	sub_wire2(212, 22)    <= sub_wire45(22);
	sub_wire2(212, 23)    <= sub_wire45(23);
	sub_wire2(212, 24)    <= sub_wire45(24);
	sub_wire2(212, 25)    <= sub_wire45(25);
	sub_wire2(212, 26)    <= sub_wire45(26);
	sub_wire2(212, 27)    <= sub_wire45(27);
	sub_wire2(212, 28)    <= sub_wire45(28);
	sub_wire2(212, 29)    <= sub_wire45(29);
	sub_wire2(212, 30)    <= sub_wire45(30);
	sub_wire2(212, 31)    <= sub_wire45(31);
	sub_wire2(212, 32)    <= sub_wire45(32);
	sub_wire2(212, 33)    <= sub_wire45(33);
	sub_wire2(212, 34)    <= sub_wire45(34);
	sub_wire2(212, 35)    <= sub_wire45(35);
	sub_wire2(212, 36)    <= sub_wire45(36);
	sub_wire2(212, 37)    <= sub_wire45(37);
	sub_wire2(212, 38)    <= sub_wire45(38);
	sub_wire2(212, 39)    <= sub_wire45(39);
	sub_wire2(211, 0)    <= sub_wire46(0);
	sub_wire2(211, 1)    <= sub_wire46(1);
	sub_wire2(211, 2)    <= sub_wire46(2);
	sub_wire2(211, 3)    <= sub_wire46(3);
	sub_wire2(211, 4)    <= sub_wire46(4);
	sub_wire2(211, 5)    <= sub_wire46(5);
	sub_wire2(211, 6)    <= sub_wire46(6);
	sub_wire2(211, 7)    <= sub_wire46(7);
	sub_wire2(211, 8)    <= sub_wire46(8);
	sub_wire2(211, 9)    <= sub_wire46(9);
	sub_wire2(211, 10)    <= sub_wire46(10);
	sub_wire2(211, 11)    <= sub_wire46(11);
	sub_wire2(211, 12)    <= sub_wire46(12);
	sub_wire2(211, 13)    <= sub_wire46(13);
	sub_wire2(211, 14)    <= sub_wire46(14);
	sub_wire2(211, 15)    <= sub_wire46(15);
	sub_wire2(211, 16)    <= sub_wire46(16);
	sub_wire2(211, 17)    <= sub_wire46(17);
	sub_wire2(211, 18)    <= sub_wire46(18);
	sub_wire2(211, 19)    <= sub_wire46(19);
	sub_wire2(211, 20)    <= sub_wire46(20);
	sub_wire2(211, 21)    <= sub_wire46(21);
	sub_wire2(211, 22)    <= sub_wire46(22);
	sub_wire2(211, 23)    <= sub_wire46(23);
	sub_wire2(211, 24)    <= sub_wire46(24);
	sub_wire2(211, 25)    <= sub_wire46(25);
	sub_wire2(211, 26)    <= sub_wire46(26);
	sub_wire2(211, 27)    <= sub_wire46(27);
	sub_wire2(211, 28)    <= sub_wire46(28);
	sub_wire2(211, 29)    <= sub_wire46(29);
	sub_wire2(211, 30)    <= sub_wire46(30);
	sub_wire2(211, 31)    <= sub_wire46(31);
	sub_wire2(211, 32)    <= sub_wire46(32);
	sub_wire2(211, 33)    <= sub_wire46(33);
	sub_wire2(211, 34)    <= sub_wire46(34);
	sub_wire2(211, 35)    <= sub_wire46(35);
	sub_wire2(211, 36)    <= sub_wire46(36);
	sub_wire2(211, 37)    <= sub_wire46(37);
	sub_wire2(211, 38)    <= sub_wire46(38);
	sub_wire2(211, 39)    <= sub_wire46(39);
	sub_wire2(210, 0)    <= sub_wire47(0);
	sub_wire2(210, 1)    <= sub_wire47(1);
	sub_wire2(210, 2)    <= sub_wire47(2);
	sub_wire2(210, 3)    <= sub_wire47(3);
	sub_wire2(210, 4)    <= sub_wire47(4);
	sub_wire2(210, 5)    <= sub_wire47(5);
	sub_wire2(210, 6)    <= sub_wire47(6);
	sub_wire2(210, 7)    <= sub_wire47(7);
	sub_wire2(210, 8)    <= sub_wire47(8);
	sub_wire2(210, 9)    <= sub_wire47(9);
	sub_wire2(210, 10)    <= sub_wire47(10);
	sub_wire2(210, 11)    <= sub_wire47(11);
	sub_wire2(210, 12)    <= sub_wire47(12);
	sub_wire2(210, 13)    <= sub_wire47(13);
	sub_wire2(210, 14)    <= sub_wire47(14);
	sub_wire2(210, 15)    <= sub_wire47(15);
	sub_wire2(210, 16)    <= sub_wire47(16);
	sub_wire2(210, 17)    <= sub_wire47(17);
	sub_wire2(210, 18)    <= sub_wire47(18);
	sub_wire2(210, 19)    <= sub_wire47(19);
	sub_wire2(210, 20)    <= sub_wire47(20);
	sub_wire2(210, 21)    <= sub_wire47(21);
	sub_wire2(210, 22)    <= sub_wire47(22);
	sub_wire2(210, 23)    <= sub_wire47(23);
	sub_wire2(210, 24)    <= sub_wire47(24);
	sub_wire2(210, 25)    <= sub_wire47(25);
	sub_wire2(210, 26)    <= sub_wire47(26);
	sub_wire2(210, 27)    <= sub_wire47(27);
	sub_wire2(210, 28)    <= sub_wire47(28);
	sub_wire2(210, 29)    <= sub_wire47(29);
	sub_wire2(210, 30)    <= sub_wire47(30);
	sub_wire2(210, 31)    <= sub_wire47(31);
	sub_wire2(210, 32)    <= sub_wire47(32);
	sub_wire2(210, 33)    <= sub_wire47(33);
	sub_wire2(210, 34)    <= sub_wire47(34);
	sub_wire2(210, 35)    <= sub_wire47(35);
	sub_wire2(210, 36)    <= sub_wire47(36);
	sub_wire2(210, 37)    <= sub_wire47(37);
	sub_wire2(210, 38)    <= sub_wire47(38);
	sub_wire2(210, 39)    <= sub_wire47(39);
	sub_wire2(209, 0)    <= sub_wire48(0);
	sub_wire2(209, 1)    <= sub_wire48(1);
	sub_wire2(209, 2)    <= sub_wire48(2);
	sub_wire2(209, 3)    <= sub_wire48(3);
	sub_wire2(209, 4)    <= sub_wire48(4);
	sub_wire2(209, 5)    <= sub_wire48(5);
	sub_wire2(209, 6)    <= sub_wire48(6);
	sub_wire2(209, 7)    <= sub_wire48(7);
	sub_wire2(209, 8)    <= sub_wire48(8);
	sub_wire2(209, 9)    <= sub_wire48(9);
	sub_wire2(209, 10)    <= sub_wire48(10);
	sub_wire2(209, 11)    <= sub_wire48(11);
	sub_wire2(209, 12)    <= sub_wire48(12);
	sub_wire2(209, 13)    <= sub_wire48(13);
	sub_wire2(209, 14)    <= sub_wire48(14);
	sub_wire2(209, 15)    <= sub_wire48(15);
	sub_wire2(209, 16)    <= sub_wire48(16);
	sub_wire2(209, 17)    <= sub_wire48(17);
	sub_wire2(209, 18)    <= sub_wire48(18);
	sub_wire2(209, 19)    <= sub_wire48(19);
	sub_wire2(209, 20)    <= sub_wire48(20);
	sub_wire2(209, 21)    <= sub_wire48(21);
	sub_wire2(209, 22)    <= sub_wire48(22);
	sub_wire2(209, 23)    <= sub_wire48(23);
	sub_wire2(209, 24)    <= sub_wire48(24);
	sub_wire2(209, 25)    <= sub_wire48(25);
	sub_wire2(209, 26)    <= sub_wire48(26);
	sub_wire2(209, 27)    <= sub_wire48(27);
	sub_wire2(209, 28)    <= sub_wire48(28);
	sub_wire2(209, 29)    <= sub_wire48(29);
	sub_wire2(209, 30)    <= sub_wire48(30);
	sub_wire2(209, 31)    <= sub_wire48(31);
	sub_wire2(209, 32)    <= sub_wire48(32);
	sub_wire2(209, 33)    <= sub_wire48(33);
	sub_wire2(209, 34)    <= sub_wire48(34);
	sub_wire2(209, 35)    <= sub_wire48(35);
	sub_wire2(209, 36)    <= sub_wire48(36);
	sub_wire2(209, 37)    <= sub_wire48(37);
	sub_wire2(209, 38)    <= sub_wire48(38);
	sub_wire2(209, 39)    <= sub_wire48(39);
	sub_wire2(208, 0)    <= sub_wire49(0);
	sub_wire2(208, 1)    <= sub_wire49(1);
	sub_wire2(208, 2)    <= sub_wire49(2);
	sub_wire2(208, 3)    <= sub_wire49(3);
	sub_wire2(208, 4)    <= sub_wire49(4);
	sub_wire2(208, 5)    <= sub_wire49(5);
	sub_wire2(208, 6)    <= sub_wire49(6);
	sub_wire2(208, 7)    <= sub_wire49(7);
	sub_wire2(208, 8)    <= sub_wire49(8);
	sub_wire2(208, 9)    <= sub_wire49(9);
	sub_wire2(208, 10)    <= sub_wire49(10);
	sub_wire2(208, 11)    <= sub_wire49(11);
	sub_wire2(208, 12)    <= sub_wire49(12);
	sub_wire2(208, 13)    <= sub_wire49(13);
	sub_wire2(208, 14)    <= sub_wire49(14);
	sub_wire2(208, 15)    <= sub_wire49(15);
	sub_wire2(208, 16)    <= sub_wire49(16);
	sub_wire2(208, 17)    <= sub_wire49(17);
	sub_wire2(208, 18)    <= sub_wire49(18);
	sub_wire2(208, 19)    <= sub_wire49(19);
	sub_wire2(208, 20)    <= sub_wire49(20);
	sub_wire2(208, 21)    <= sub_wire49(21);
	sub_wire2(208, 22)    <= sub_wire49(22);
	sub_wire2(208, 23)    <= sub_wire49(23);
	sub_wire2(208, 24)    <= sub_wire49(24);
	sub_wire2(208, 25)    <= sub_wire49(25);
	sub_wire2(208, 26)    <= sub_wire49(26);
	sub_wire2(208, 27)    <= sub_wire49(27);
	sub_wire2(208, 28)    <= sub_wire49(28);
	sub_wire2(208, 29)    <= sub_wire49(29);
	sub_wire2(208, 30)    <= sub_wire49(30);
	sub_wire2(208, 31)    <= sub_wire49(31);
	sub_wire2(208, 32)    <= sub_wire49(32);
	sub_wire2(208, 33)    <= sub_wire49(33);
	sub_wire2(208, 34)    <= sub_wire49(34);
	sub_wire2(208, 35)    <= sub_wire49(35);
	sub_wire2(208, 36)    <= sub_wire49(36);
	sub_wire2(208, 37)    <= sub_wire49(37);
	sub_wire2(208, 38)    <= sub_wire49(38);
	sub_wire2(208, 39)    <= sub_wire49(39);
	sub_wire2(207, 0)    <= sub_wire50(0);
	sub_wire2(207, 1)    <= sub_wire50(1);
	sub_wire2(207, 2)    <= sub_wire50(2);
	sub_wire2(207, 3)    <= sub_wire50(3);
	sub_wire2(207, 4)    <= sub_wire50(4);
	sub_wire2(207, 5)    <= sub_wire50(5);
	sub_wire2(207, 6)    <= sub_wire50(6);
	sub_wire2(207, 7)    <= sub_wire50(7);
	sub_wire2(207, 8)    <= sub_wire50(8);
	sub_wire2(207, 9)    <= sub_wire50(9);
	sub_wire2(207, 10)    <= sub_wire50(10);
	sub_wire2(207, 11)    <= sub_wire50(11);
	sub_wire2(207, 12)    <= sub_wire50(12);
	sub_wire2(207, 13)    <= sub_wire50(13);
	sub_wire2(207, 14)    <= sub_wire50(14);
	sub_wire2(207, 15)    <= sub_wire50(15);
	sub_wire2(207, 16)    <= sub_wire50(16);
	sub_wire2(207, 17)    <= sub_wire50(17);
	sub_wire2(207, 18)    <= sub_wire50(18);
	sub_wire2(207, 19)    <= sub_wire50(19);
	sub_wire2(207, 20)    <= sub_wire50(20);
	sub_wire2(207, 21)    <= sub_wire50(21);
	sub_wire2(207, 22)    <= sub_wire50(22);
	sub_wire2(207, 23)    <= sub_wire50(23);
	sub_wire2(207, 24)    <= sub_wire50(24);
	sub_wire2(207, 25)    <= sub_wire50(25);
	sub_wire2(207, 26)    <= sub_wire50(26);
	sub_wire2(207, 27)    <= sub_wire50(27);
	sub_wire2(207, 28)    <= sub_wire50(28);
	sub_wire2(207, 29)    <= sub_wire50(29);
	sub_wire2(207, 30)    <= sub_wire50(30);
	sub_wire2(207, 31)    <= sub_wire50(31);
	sub_wire2(207, 32)    <= sub_wire50(32);
	sub_wire2(207, 33)    <= sub_wire50(33);
	sub_wire2(207, 34)    <= sub_wire50(34);
	sub_wire2(207, 35)    <= sub_wire50(35);
	sub_wire2(207, 36)    <= sub_wire50(36);
	sub_wire2(207, 37)    <= sub_wire50(37);
	sub_wire2(207, 38)    <= sub_wire50(38);
	sub_wire2(207, 39)    <= sub_wire50(39);
	sub_wire2(206, 0)    <= sub_wire51(0);
	sub_wire2(206, 1)    <= sub_wire51(1);
	sub_wire2(206, 2)    <= sub_wire51(2);
	sub_wire2(206, 3)    <= sub_wire51(3);
	sub_wire2(206, 4)    <= sub_wire51(4);
	sub_wire2(206, 5)    <= sub_wire51(5);
	sub_wire2(206, 6)    <= sub_wire51(6);
	sub_wire2(206, 7)    <= sub_wire51(7);
	sub_wire2(206, 8)    <= sub_wire51(8);
	sub_wire2(206, 9)    <= sub_wire51(9);
	sub_wire2(206, 10)    <= sub_wire51(10);
	sub_wire2(206, 11)    <= sub_wire51(11);
	sub_wire2(206, 12)    <= sub_wire51(12);
	sub_wire2(206, 13)    <= sub_wire51(13);
	sub_wire2(206, 14)    <= sub_wire51(14);
	sub_wire2(206, 15)    <= sub_wire51(15);
	sub_wire2(206, 16)    <= sub_wire51(16);
	sub_wire2(206, 17)    <= sub_wire51(17);
	sub_wire2(206, 18)    <= sub_wire51(18);
	sub_wire2(206, 19)    <= sub_wire51(19);
	sub_wire2(206, 20)    <= sub_wire51(20);
	sub_wire2(206, 21)    <= sub_wire51(21);
	sub_wire2(206, 22)    <= sub_wire51(22);
	sub_wire2(206, 23)    <= sub_wire51(23);
	sub_wire2(206, 24)    <= sub_wire51(24);
	sub_wire2(206, 25)    <= sub_wire51(25);
	sub_wire2(206, 26)    <= sub_wire51(26);
	sub_wire2(206, 27)    <= sub_wire51(27);
	sub_wire2(206, 28)    <= sub_wire51(28);
	sub_wire2(206, 29)    <= sub_wire51(29);
	sub_wire2(206, 30)    <= sub_wire51(30);
	sub_wire2(206, 31)    <= sub_wire51(31);
	sub_wire2(206, 32)    <= sub_wire51(32);
	sub_wire2(206, 33)    <= sub_wire51(33);
	sub_wire2(206, 34)    <= sub_wire51(34);
	sub_wire2(206, 35)    <= sub_wire51(35);
	sub_wire2(206, 36)    <= sub_wire51(36);
	sub_wire2(206, 37)    <= sub_wire51(37);
	sub_wire2(206, 38)    <= sub_wire51(38);
	sub_wire2(206, 39)    <= sub_wire51(39);
	sub_wire2(205, 0)    <= sub_wire52(0);
	sub_wire2(205, 1)    <= sub_wire52(1);
	sub_wire2(205, 2)    <= sub_wire52(2);
	sub_wire2(205, 3)    <= sub_wire52(3);
	sub_wire2(205, 4)    <= sub_wire52(4);
	sub_wire2(205, 5)    <= sub_wire52(5);
	sub_wire2(205, 6)    <= sub_wire52(6);
	sub_wire2(205, 7)    <= sub_wire52(7);
	sub_wire2(205, 8)    <= sub_wire52(8);
	sub_wire2(205, 9)    <= sub_wire52(9);
	sub_wire2(205, 10)    <= sub_wire52(10);
	sub_wire2(205, 11)    <= sub_wire52(11);
	sub_wire2(205, 12)    <= sub_wire52(12);
	sub_wire2(205, 13)    <= sub_wire52(13);
	sub_wire2(205, 14)    <= sub_wire52(14);
	sub_wire2(205, 15)    <= sub_wire52(15);
	sub_wire2(205, 16)    <= sub_wire52(16);
	sub_wire2(205, 17)    <= sub_wire52(17);
	sub_wire2(205, 18)    <= sub_wire52(18);
	sub_wire2(205, 19)    <= sub_wire52(19);
	sub_wire2(205, 20)    <= sub_wire52(20);
	sub_wire2(205, 21)    <= sub_wire52(21);
	sub_wire2(205, 22)    <= sub_wire52(22);
	sub_wire2(205, 23)    <= sub_wire52(23);
	sub_wire2(205, 24)    <= sub_wire52(24);
	sub_wire2(205, 25)    <= sub_wire52(25);
	sub_wire2(205, 26)    <= sub_wire52(26);
	sub_wire2(205, 27)    <= sub_wire52(27);
	sub_wire2(205, 28)    <= sub_wire52(28);
	sub_wire2(205, 29)    <= sub_wire52(29);
	sub_wire2(205, 30)    <= sub_wire52(30);
	sub_wire2(205, 31)    <= sub_wire52(31);
	sub_wire2(205, 32)    <= sub_wire52(32);
	sub_wire2(205, 33)    <= sub_wire52(33);
	sub_wire2(205, 34)    <= sub_wire52(34);
	sub_wire2(205, 35)    <= sub_wire52(35);
	sub_wire2(205, 36)    <= sub_wire52(36);
	sub_wire2(205, 37)    <= sub_wire52(37);
	sub_wire2(205, 38)    <= sub_wire52(38);
	sub_wire2(205, 39)    <= sub_wire52(39);
	sub_wire2(204, 0)    <= sub_wire53(0);
	sub_wire2(204, 1)    <= sub_wire53(1);
	sub_wire2(204, 2)    <= sub_wire53(2);
	sub_wire2(204, 3)    <= sub_wire53(3);
	sub_wire2(204, 4)    <= sub_wire53(4);
	sub_wire2(204, 5)    <= sub_wire53(5);
	sub_wire2(204, 6)    <= sub_wire53(6);
	sub_wire2(204, 7)    <= sub_wire53(7);
	sub_wire2(204, 8)    <= sub_wire53(8);
	sub_wire2(204, 9)    <= sub_wire53(9);
	sub_wire2(204, 10)    <= sub_wire53(10);
	sub_wire2(204, 11)    <= sub_wire53(11);
	sub_wire2(204, 12)    <= sub_wire53(12);
	sub_wire2(204, 13)    <= sub_wire53(13);
	sub_wire2(204, 14)    <= sub_wire53(14);
	sub_wire2(204, 15)    <= sub_wire53(15);
	sub_wire2(204, 16)    <= sub_wire53(16);
	sub_wire2(204, 17)    <= sub_wire53(17);
	sub_wire2(204, 18)    <= sub_wire53(18);
	sub_wire2(204, 19)    <= sub_wire53(19);
	sub_wire2(204, 20)    <= sub_wire53(20);
	sub_wire2(204, 21)    <= sub_wire53(21);
	sub_wire2(204, 22)    <= sub_wire53(22);
	sub_wire2(204, 23)    <= sub_wire53(23);
	sub_wire2(204, 24)    <= sub_wire53(24);
	sub_wire2(204, 25)    <= sub_wire53(25);
	sub_wire2(204, 26)    <= sub_wire53(26);
	sub_wire2(204, 27)    <= sub_wire53(27);
	sub_wire2(204, 28)    <= sub_wire53(28);
	sub_wire2(204, 29)    <= sub_wire53(29);
	sub_wire2(204, 30)    <= sub_wire53(30);
	sub_wire2(204, 31)    <= sub_wire53(31);
	sub_wire2(204, 32)    <= sub_wire53(32);
	sub_wire2(204, 33)    <= sub_wire53(33);
	sub_wire2(204, 34)    <= sub_wire53(34);
	sub_wire2(204, 35)    <= sub_wire53(35);
	sub_wire2(204, 36)    <= sub_wire53(36);
	sub_wire2(204, 37)    <= sub_wire53(37);
	sub_wire2(204, 38)    <= sub_wire53(38);
	sub_wire2(204, 39)    <= sub_wire53(39);
	sub_wire2(203, 0)    <= sub_wire54(0);
	sub_wire2(203, 1)    <= sub_wire54(1);
	sub_wire2(203, 2)    <= sub_wire54(2);
	sub_wire2(203, 3)    <= sub_wire54(3);
	sub_wire2(203, 4)    <= sub_wire54(4);
	sub_wire2(203, 5)    <= sub_wire54(5);
	sub_wire2(203, 6)    <= sub_wire54(6);
	sub_wire2(203, 7)    <= sub_wire54(7);
	sub_wire2(203, 8)    <= sub_wire54(8);
	sub_wire2(203, 9)    <= sub_wire54(9);
	sub_wire2(203, 10)    <= sub_wire54(10);
	sub_wire2(203, 11)    <= sub_wire54(11);
	sub_wire2(203, 12)    <= sub_wire54(12);
	sub_wire2(203, 13)    <= sub_wire54(13);
	sub_wire2(203, 14)    <= sub_wire54(14);
	sub_wire2(203, 15)    <= sub_wire54(15);
	sub_wire2(203, 16)    <= sub_wire54(16);
	sub_wire2(203, 17)    <= sub_wire54(17);
	sub_wire2(203, 18)    <= sub_wire54(18);
	sub_wire2(203, 19)    <= sub_wire54(19);
	sub_wire2(203, 20)    <= sub_wire54(20);
	sub_wire2(203, 21)    <= sub_wire54(21);
	sub_wire2(203, 22)    <= sub_wire54(22);
	sub_wire2(203, 23)    <= sub_wire54(23);
	sub_wire2(203, 24)    <= sub_wire54(24);
	sub_wire2(203, 25)    <= sub_wire54(25);
	sub_wire2(203, 26)    <= sub_wire54(26);
	sub_wire2(203, 27)    <= sub_wire54(27);
	sub_wire2(203, 28)    <= sub_wire54(28);
	sub_wire2(203, 29)    <= sub_wire54(29);
	sub_wire2(203, 30)    <= sub_wire54(30);
	sub_wire2(203, 31)    <= sub_wire54(31);
	sub_wire2(203, 32)    <= sub_wire54(32);
	sub_wire2(203, 33)    <= sub_wire54(33);
	sub_wire2(203, 34)    <= sub_wire54(34);
	sub_wire2(203, 35)    <= sub_wire54(35);
	sub_wire2(203, 36)    <= sub_wire54(36);
	sub_wire2(203, 37)    <= sub_wire54(37);
	sub_wire2(203, 38)    <= sub_wire54(38);
	sub_wire2(203, 39)    <= sub_wire54(39);
	sub_wire2(202, 0)    <= sub_wire55(0);
	sub_wire2(202, 1)    <= sub_wire55(1);
	sub_wire2(202, 2)    <= sub_wire55(2);
	sub_wire2(202, 3)    <= sub_wire55(3);
	sub_wire2(202, 4)    <= sub_wire55(4);
	sub_wire2(202, 5)    <= sub_wire55(5);
	sub_wire2(202, 6)    <= sub_wire55(6);
	sub_wire2(202, 7)    <= sub_wire55(7);
	sub_wire2(202, 8)    <= sub_wire55(8);
	sub_wire2(202, 9)    <= sub_wire55(9);
	sub_wire2(202, 10)    <= sub_wire55(10);
	sub_wire2(202, 11)    <= sub_wire55(11);
	sub_wire2(202, 12)    <= sub_wire55(12);
	sub_wire2(202, 13)    <= sub_wire55(13);
	sub_wire2(202, 14)    <= sub_wire55(14);
	sub_wire2(202, 15)    <= sub_wire55(15);
	sub_wire2(202, 16)    <= sub_wire55(16);
	sub_wire2(202, 17)    <= sub_wire55(17);
	sub_wire2(202, 18)    <= sub_wire55(18);
	sub_wire2(202, 19)    <= sub_wire55(19);
	sub_wire2(202, 20)    <= sub_wire55(20);
	sub_wire2(202, 21)    <= sub_wire55(21);
	sub_wire2(202, 22)    <= sub_wire55(22);
	sub_wire2(202, 23)    <= sub_wire55(23);
	sub_wire2(202, 24)    <= sub_wire55(24);
	sub_wire2(202, 25)    <= sub_wire55(25);
	sub_wire2(202, 26)    <= sub_wire55(26);
	sub_wire2(202, 27)    <= sub_wire55(27);
	sub_wire2(202, 28)    <= sub_wire55(28);
	sub_wire2(202, 29)    <= sub_wire55(29);
	sub_wire2(202, 30)    <= sub_wire55(30);
	sub_wire2(202, 31)    <= sub_wire55(31);
	sub_wire2(202, 32)    <= sub_wire55(32);
	sub_wire2(202, 33)    <= sub_wire55(33);
	sub_wire2(202, 34)    <= sub_wire55(34);
	sub_wire2(202, 35)    <= sub_wire55(35);
	sub_wire2(202, 36)    <= sub_wire55(36);
	sub_wire2(202, 37)    <= sub_wire55(37);
	sub_wire2(202, 38)    <= sub_wire55(38);
	sub_wire2(202, 39)    <= sub_wire55(39);
	sub_wire2(201, 0)    <= sub_wire56(0);
	sub_wire2(201, 1)    <= sub_wire56(1);
	sub_wire2(201, 2)    <= sub_wire56(2);
	sub_wire2(201, 3)    <= sub_wire56(3);
	sub_wire2(201, 4)    <= sub_wire56(4);
	sub_wire2(201, 5)    <= sub_wire56(5);
	sub_wire2(201, 6)    <= sub_wire56(6);
	sub_wire2(201, 7)    <= sub_wire56(7);
	sub_wire2(201, 8)    <= sub_wire56(8);
	sub_wire2(201, 9)    <= sub_wire56(9);
	sub_wire2(201, 10)    <= sub_wire56(10);
	sub_wire2(201, 11)    <= sub_wire56(11);
	sub_wire2(201, 12)    <= sub_wire56(12);
	sub_wire2(201, 13)    <= sub_wire56(13);
	sub_wire2(201, 14)    <= sub_wire56(14);
	sub_wire2(201, 15)    <= sub_wire56(15);
	sub_wire2(201, 16)    <= sub_wire56(16);
	sub_wire2(201, 17)    <= sub_wire56(17);
	sub_wire2(201, 18)    <= sub_wire56(18);
	sub_wire2(201, 19)    <= sub_wire56(19);
	sub_wire2(201, 20)    <= sub_wire56(20);
	sub_wire2(201, 21)    <= sub_wire56(21);
	sub_wire2(201, 22)    <= sub_wire56(22);
	sub_wire2(201, 23)    <= sub_wire56(23);
	sub_wire2(201, 24)    <= sub_wire56(24);
	sub_wire2(201, 25)    <= sub_wire56(25);
	sub_wire2(201, 26)    <= sub_wire56(26);
	sub_wire2(201, 27)    <= sub_wire56(27);
	sub_wire2(201, 28)    <= sub_wire56(28);
	sub_wire2(201, 29)    <= sub_wire56(29);
	sub_wire2(201, 30)    <= sub_wire56(30);
	sub_wire2(201, 31)    <= sub_wire56(31);
	sub_wire2(201, 32)    <= sub_wire56(32);
	sub_wire2(201, 33)    <= sub_wire56(33);
	sub_wire2(201, 34)    <= sub_wire56(34);
	sub_wire2(201, 35)    <= sub_wire56(35);
	sub_wire2(201, 36)    <= sub_wire56(36);
	sub_wire2(201, 37)    <= sub_wire56(37);
	sub_wire2(201, 38)    <= sub_wire56(38);
	sub_wire2(201, 39)    <= sub_wire56(39);
	sub_wire2(200, 0)    <= sub_wire57(0);
	sub_wire2(200, 1)    <= sub_wire57(1);
	sub_wire2(200, 2)    <= sub_wire57(2);
	sub_wire2(200, 3)    <= sub_wire57(3);
	sub_wire2(200, 4)    <= sub_wire57(4);
	sub_wire2(200, 5)    <= sub_wire57(5);
	sub_wire2(200, 6)    <= sub_wire57(6);
	sub_wire2(200, 7)    <= sub_wire57(7);
	sub_wire2(200, 8)    <= sub_wire57(8);
	sub_wire2(200, 9)    <= sub_wire57(9);
	sub_wire2(200, 10)    <= sub_wire57(10);
	sub_wire2(200, 11)    <= sub_wire57(11);
	sub_wire2(200, 12)    <= sub_wire57(12);
	sub_wire2(200, 13)    <= sub_wire57(13);
	sub_wire2(200, 14)    <= sub_wire57(14);
	sub_wire2(200, 15)    <= sub_wire57(15);
	sub_wire2(200, 16)    <= sub_wire57(16);
	sub_wire2(200, 17)    <= sub_wire57(17);
	sub_wire2(200, 18)    <= sub_wire57(18);
	sub_wire2(200, 19)    <= sub_wire57(19);
	sub_wire2(200, 20)    <= sub_wire57(20);
	sub_wire2(200, 21)    <= sub_wire57(21);
	sub_wire2(200, 22)    <= sub_wire57(22);
	sub_wire2(200, 23)    <= sub_wire57(23);
	sub_wire2(200, 24)    <= sub_wire57(24);
	sub_wire2(200, 25)    <= sub_wire57(25);
	sub_wire2(200, 26)    <= sub_wire57(26);
	sub_wire2(200, 27)    <= sub_wire57(27);
	sub_wire2(200, 28)    <= sub_wire57(28);
	sub_wire2(200, 29)    <= sub_wire57(29);
	sub_wire2(200, 30)    <= sub_wire57(30);
	sub_wire2(200, 31)    <= sub_wire57(31);
	sub_wire2(200, 32)    <= sub_wire57(32);
	sub_wire2(200, 33)    <= sub_wire57(33);
	sub_wire2(200, 34)    <= sub_wire57(34);
	sub_wire2(200, 35)    <= sub_wire57(35);
	sub_wire2(200, 36)    <= sub_wire57(36);
	sub_wire2(200, 37)    <= sub_wire57(37);
	sub_wire2(200, 38)    <= sub_wire57(38);
	sub_wire2(200, 39)    <= sub_wire57(39);
	sub_wire2(199, 0)    <= sub_wire58(0);
	sub_wire2(199, 1)    <= sub_wire58(1);
	sub_wire2(199, 2)    <= sub_wire58(2);
	sub_wire2(199, 3)    <= sub_wire58(3);
	sub_wire2(199, 4)    <= sub_wire58(4);
	sub_wire2(199, 5)    <= sub_wire58(5);
	sub_wire2(199, 6)    <= sub_wire58(6);
	sub_wire2(199, 7)    <= sub_wire58(7);
	sub_wire2(199, 8)    <= sub_wire58(8);
	sub_wire2(199, 9)    <= sub_wire58(9);
	sub_wire2(199, 10)    <= sub_wire58(10);
	sub_wire2(199, 11)    <= sub_wire58(11);
	sub_wire2(199, 12)    <= sub_wire58(12);
	sub_wire2(199, 13)    <= sub_wire58(13);
	sub_wire2(199, 14)    <= sub_wire58(14);
	sub_wire2(199, 15)    <= sub_wire58(15);
	sub_wire2(199, 16)    <= sub_wire58(16);
	sub_wire2(199, 17)    <= sub_wire58(17);
	sub_wire2(199, 18)    <= sub_wire58(18);
	sub_wire2(199, 19)    <= sub_wire58(19);
	sub_wire2(199, 20)    <= sub_wire58(20);
	sub_wire2(199, 21)    <= sub_wire58(21);
	sub_wire2(199, 22)    <= sub_wire58(22);
	sub_wire2(199, 23)    <= sub_wire58(23);
	sub_wire2(199, 24)    <= sub_wire58(24);
	sub_wire2(199, 25)    <= sub_wire58(25);
	sub_wire2(199, 26)    <= sub_wire58(26);
	sub_wire2(199, 27)    <= sub_wire58(27);
	sub_wire2(199, 28)    <= sub_wire58(28);
	sub_wire2(199, 29)    <= sub_wire58(29);
	sub_wire2(199, 30)    <= sub_wire58(30);
	sub_wire2(199, 31)    <= sub_wire58(31);
	sub_wire2(199, 32)    <= sub_wire58(32);
	sub_wire2(199, 33)    <= sub_wire58(33);
	sub_wire2(199, 34)    <= sub_wire58(34);
	sub_wire2(199, 35)    <= sub_wire58(35);
	sub_wire2(199, 36)    <= sub_wire58(36);
	sub_wire2(199, 37)    <= sub_wire58(37);
	sub_wire2(199, 38)    <= sub_wire58(38);
	sub_wire2(199, 39)    <= sub_wire58(39);
	sub_wire2(198, 0)    <= sub_wire59(0);
	sub_wire2(198, 1)    <= sub_wire59(1);
	sub_wire2(198, 2)    <= sub_wire59(2);
	sub_wire2(198, 3)    <= sub_wire59(3);
	sub_wire2(198, 4)    <= sub_wire59(4);
	sub_wire2(198, 5)    <= sub_wire59(5);
	sub_wire2(198, 6)    <= sub_wire59(6);
	sub_wire2(198, 7)    <= sub_wire59(7);
	sub_wire2(198, 8)    <= sub_wire59(8);
	sub_wire2(198, 9)    <= sub_wire59(9);
	sub_wire2(198, 10)    <= sub_wire59(10);
	sub_wire2(198, 11)    <= sub_wire59(11);
	sub_wire2(198, 12)    <= sub_wire59(12);
	sub_wire2(198, 13)    <= sub_wire59(13);
	sub_wire2(198, 14)    <= sub_wire59(14);
	sub_wire2(198, 15)    <= sub_wire59(15);
	sub_wire2(198, 16)    <= sub_wire59(16);
	sub_wire2(198, 17)    <= sub_wire59(17);
	sub_wire2(198, 18)    <= sub_wire59(18);
	sub_wire2(198, 19)    <= sub_wire59(19);
	sub_wire2(198, 20)    <= sub_wire59(20);
	sub_wire2(198, 21)    <= sub_wire59(21);
	sub_wire2(198, 22)    <= sub_wire59(22);
	sub_wire2(198, 23)    <= sub_wire59(23);
	sub_wire2(198, 24)    <= sub_wire59(24);
	sub_wire2(198, 25)    <= sub_wire59(25);
	sub_wire2(198, 26)    <= sub_wire59(26);
	sub_wire2(198, 27)    <= sub_wire59(27);
	sub_wire2(198, 28)    <= sub_wire59(28);
	sub_wire2(198, 29)    <= sub_wire59(29);
	sub_wire2(198, 30)    <= sub_wire59(30);
	sub_wire2(198, 31)    <= sub_wire59(31);
	sub_wire2(198, 32)    <= sub_wire59(32);
	sub_wire2(198, 33)    <= sub_wire59(33);
	sub_wire2(198, 34)    <= sub_wire59(34);
	sub_wire2(198, 35)    <= sub_wire59(35);
	sub_wire2(198, 36)    <= sub_wire59(36);
	sub_wire2(198, 37)    <= sub_wire59(37);
	sub_wire2(198, 38)    <= sub_wire59(38);
	sub_wire2(198, 39)    <= sub_wire59(39);
	sub_wire2(197, 0)    <= sub_wire60(0);
	sub_wire2(197, 1)    <= sub_wire60(1);
	sub_wire2(197, 2)    <= sub_wire60(2);
	sub_wire2(197, 3)    <= sub_wire60(3);
	sub_wire2(197, 4)    <= sub_wire60(4);
	sub_wire2(197, 5)    <= sub_wire60(5);
	sub_wire2(197, 6)    <= sub_wire60(6);
	sub_wire2(197, 7)    <= sub_wire60(7);
	sub_wire2(197, 8)    <= sub_wire60(8);
	sub_wire2(197, 9)    <= sub_wire60(9);
	sub_wire2(197, 10)    <= sub_wire60(10);
	sub_wire2(197, 11)    <= sub_wire60(11);
	sub_wire2(197, 12)    <= sub_wire60(12);
	sub_wire2(197, 13)    <= sub_wire60(13);
	sub_wire2(197, 14)    <= sub_wire60(14);
	sub_wire2(197, 15)    <= sub_wire60(15);
	sub_wire2(197, 16)    <= sub_wire60(16);
	sub_wire2(197, 17)    <= sub_wire60(17);
	sub_wire2(197, 18)    <= sub_wire60(18);
	sub_wire2(197, 19)    <= sub_wire60(19);
	sub_wire2(197, 20)    <= sub_wire60(20);
	sub_wire2(197, 21)    <= sub_wire60(21);
	sub_wire2(197, 22)    <= sub_wire60(22);
	sub_wire2(197, 23)    <= sub_wire60(23);
	sub_wire2(197, 24)    <= sub_wire60(24);
	sub_wire2(197, 25)    <= sub_wire60(25);
	sub_wire2(197, 26)    <= sub_wire60(26);
	sub_wire2(197, 27)    <= sub_wire60(27);
	sub_wire2(197, 28)    <= sub_wire60(28);
	sub_wire2(197, 29)    <= sub_wire60(29);
	sub_wire2(197, 30)    <= sub_wire60(30);
	sub_wire2(197, 31)    <= sub_wire60(31);
	sub_wire2(197, 32)    <= sub_wire60(32);
	sub_wire2(197, 33)    <= sub_wire60(33);
	sub_wire2(197, 34)    <= sub_wire60(34);
	sub_wire2(197, 35)    <= sub_wire60(35);
	sub_wire2(197, 36)    <= sub_wire60(36);
	sub_wire2(197, 37)    <= sub_wire60(37);
	sub_wire2(197, 38)    <= sub_wire60(38);
	sub_wire2(197, 39)    <= sub_wire60(39);
	sub_wire2(196, 0)    <= sub_wire61(0);
	sub_wire2(196, 1)    <= sub_wire61(1);
	sub_wire2(196, 2)    <= sub_wire61(2);
	sub_wire2(196, 3)    <= sub_wire61(3);
	sub_wire2(196, 4)    <= sub_wire61(4);
	sub_wire2(196, 5)    <= sub_wire61(5);
	sub_wire2(196, 6)    <= sub_wire61(6);
	sub_wire2(196, 7)    <= sub_wire61(7);
	sub_wire2(196, 8)    <= sub_wire61(8);
	sub_wire2(196, 9)    <= sub_wire61(9);
	sub_wire2(196, 10)    <= sub_wire61(10);
	sub_wire2(196, 11)    <= sub_wire61(11);
	sub_wire2(196, 12)    <= sub_wire61(12);
	sub_wire2(196, 13)    <= sub_wire61(13);
	sub_wire2(196, 14)    <= sub_wire61(14);
	sub_wire2(196, 15)    <= sub_wire61(15);
	sub_wire2(196, 16)    <= sub_wire61(16);
	sub_wire2(196, 17)    <= sub_wire61(17);
	sub_wire2(196, 18)    <= sub_wire61(18);
	sub_wire2(196, 19)    <= sub_wire61(19);
	sub_wire2(196, 20)    <= sub_wire61(20);
	sub_wire2(196, 21)    <= sub_wire61(21);
	sub_wire2(196, 22)    <= sub_wire61(22);
	sub_wire2(196, 23)    <= sub_wire61(23);
	sub_wire2(196, 24)    <= sub_wire61(24);
	sub_wire2(196, 25)    <= sub_wire61(25);
	sub_wire2(196, 26)    <= sub_wire61(26);
	sub_wire2(196, 27)    <= sub_wire61(27);
	sub_wire2(196, 28)    <= sub_wire61(28);
	sub_wire2(196, 29)    <= sub_wire61(29);
	sub_wire2(196, 30)    <= sub_wire61(30);
	sub_wire2(196, 31)    <= sub_wire61(31);
	sub_wire2(196, 32)    <= sub_wire61(32);
	sub_wire2(196, 33)    <= sub_wire61(33);
	sub_wire2(196, 34)    <= sub_wire61(34);
	sub_wire2(196, 35)    <= sub_wire61(35);
	sub_wire2(196, 36)    <= sub_wire61(36);
	sub_wire2(196, 37)    <= sub_wire61(37);
	sub_wire2(196, 38)    <= sub_wire61(38);
	sub_wire2(196, 39)    <= sub_wire61(39);
	sub_wire2(195, 0)    <= sub_wire62(0);
	sub_wire2(195, 1)    <= sub_wire62(1);
	sub_wire2(195, 2)    <= sub_wire62(2);
	sub_wire2(195, 3)    <= sub_wire62(3);
	sub_wire2(195, 4)    <= sub_wire62(4);
	sub_wire2(195, 5)    <= sub_wire62(5);
	sub_wire2(195, 6)    <= sub_wire62(6);
	sub_wire2(195, 7)    <= sub_wire62(7);
	sub_wire2(195, 8)    <= sub_wire62(8);
	sub_wire2(195, 9)    <= sub_wire62(9);
	sub_wire2(195, 10)    <= sub_wire62(10);
	sub_wire2(195, 11)    <= sub_wire62(11);
	sub_wire2(195, 12)    <= sub_wire62(12);
	sub_wire2(195, 13)    <= sub_wire62(13);
	sub_wire2(195, 14)    <= sub_wire62(14);
	sub_wire2(195, 15)    <= sub_wire62(15);
	sub_wire2(195, 16)    <= sub_wire62(16);
	sub_wire2(195, 17)    <= sub_wire62(17);
	sub_wire2(195, 18)    <= sub_wire62(18);
	sub_wire2(195, 19)    <= sub_wire62(19);
	sub_wire2(195, 20)    <= sub_wire62(20);
	sub_wire2(195, 21)    <= sub_wire62(21);
	sub_wire2(195, 22)    <= sub_wire62(22);
	sub_wire2(195, 23)    <= sub_wire62(23);
	sub_wire2(195, 24)    <= sub_wire62(24);
	sub_wire2(195, 25)    <= sub_wire62(25);
	sub_wire2(195, 26)    <= sub_wire62(26);
	sub_wire2(195, 27)    <= sub_wire62(27);
	sub_wire2(195, 28)    <= sub_wire62(28);
	sub_wire2(195, 29)    <= sub_wire62(29);
	sub_wire2(195, 30)    <= sub_wire62(30);
	sub_wire2(195, 31)    <= sub_wire62(31);
	sub_wire2(195, 32)    <= sub_wire62(32);
	sub_wire2(195, 33)    <= sub_wire62(33);
	sub_wire2(195, 34)    <= sub_wire62(34);
	sub_wire2(195, 35)    <= sub_wire62(35);
	sub_wire2(195, 36)    <= sub_wire62(36);
	sub_wire2(195, 37)    <= sub_wire62(37);
	sub_wire2(195, 38)    <= sub_wire62(38);
	sub_wire2(195, 39)    <= sub_wire62(39);
	sub_wire2(194, 0)    <= sub_wire63(0);
	sub_wire2(194, 1)    <= sub_wire63(1);
	sub_wire2(194, 2)    <= sub_wire63(2);
	sub_wire2(194, 3)    <= sub_wire63(3);
	sub_wire2(194, 4)    <= sub_wire63(4);
	sub_wire2(194, 5)    <= sub_wire63(5);
	sub_wire2(194, 6)    <= sub_wire63(6);
	sub_wire2(194, 7)    <= sub_wire63(7);
	sub_wire2(194, 8)    <= sub_wire63(8);
	sub_wire2(194, 9)    <= sub_wire63(9);
	sub_wire2(194, 10)    <= sub_wire63(10);
	sub_wire2(194, 11)    <= sub_wire63(11);
	sub_wire2(194, 12)    <= sub_wire63(12);
	sub_wire2(194, 13)    <= sub_wire63(13);
	sub_wire2(194, 14)    <= sub_wire63(14);
	sub_wire2(194, 15)    <= sub_wire63(15);
	sub_wire2(194, 16)    <= sub_wire63(16);
	sub_wire2(194, 17)    <= sub_wire63(17);
	sub_wire2(194, 18)    <= sub_wire63(18);
	sub_wire2(194, 19)    <= sub_wire63(19);
	sub_wire2(194, 20)    <= sub_wire63(20);
	sub_wire2(194, 21)    <= sub_wire63(21);
	sub_wire2(194, 22)    <= sub_wire63(22);
	sub_wire2(194, 23)    <= sub_wire63(23);
	sub_wire2(194, 24)    <= sub_wire63(24);
	sub_wire2(194, 25)    <= sub_wire63(25);
	sub_wire2(194, 26)    <= sub_wire63(26);
	sub_wire2(194, 27)    <= sub_wire63(27);
	sub_wire2(194, 28)    <= sub_wire63(28);
	sub_wire2(194, 29)    <= sub_wire63(29);
	sub_wire2(194, 30)    <= sub_wire63(30);
	sub_wire2(194, 31)    <= sub_wire63(31);
	sub_wire2(194, 32)    <= sub_wire63(32);
	sub_wire2(194, 33)    <= sub_wire63(33);
	sub_wire2(194, 34)    <= sub_wire63(34);
	sub_wire2(194, 35)    <= sub_wire63(35);
	sub_wire2(194, 36)    <= sub_wire63(36);
	sub_wire2(194, 37)    <= sub_wire63(37);
	sub_wire2(194, 38)    <= sub_wire63(38);
	sub_wire2(194, 39)    <= sub_wire63(39);
	sub_wire2(193, 0)    <= sub_wire64(0);
	sub_wire2(193, 1)    <= sub_wire64(1);
	sub_wire2(193, 2)    <= sub_wire64(2);
	sub_wire2(193, 3)    <= sub_wire64(3);
	sub_wire2(193, 4)    <= sub_wire64(4);
	sub_wire2(193, 5)    <= sub_wire64(5);
	sub_wire2(193, 6)    <= sub_wire64(6);
	sub_wire2(193, 7)    <= sub_wire64(7);
	sub_wire2(193, 8)    <= sub_wire64(8);
	sub_wire2(193, 9)    <= sub_wire64(9);
	sub_wire2(193, 10)    <= sub_wire64(10);
	sub_wire2(193, 11)    <= sub_wire64(11);
	sub_wire2(193, 12)    <= sub_wire64(12);
	sub_wire2(193, 13)    <= sub_wire64(13);
	sub_wire2(193, 14)    <= sub_wire64(14);
	sub_wire2(193, 15)    <= sub_wire64(15);
	sub_wire2(193, 16)    <= sub_wire64(16);
	sub_wire2(193, 17)    <= sub_wire64(17);
	sub_wire2(193, 18)    <= sub_wire64(18);
	sub_wire2(193, 19)    <= sub_wire64(19);
	sub_wire2(193, 20)    <= sub_wire64(20);
	sub_wire2(193, 21)    <= sub_wire64(21);
	sub_wire2(193, 22)    <= sub_wire64(22);
	sub_wire2(193, 23)    <= sub_wire64(23);
	sub_wire2(193, 24)    <= sub_wire64(24);
	sub_wire2(193, 25)    <= sub_wire64(25);
	sub_wire2(193, 26)    <= sub_wire64(26);
	sub_wire2(193, 27)    <= sub_wire64(27);
	sub_wire2(193, 28)    <= sub_wire64(28);
	sub_wire2(193, 29)    <= sub_wire64(29);
	sub_wire2(193, 30)    <= sub_wire64(30);
	sub_wire2(193, 31)    <= sub_wire64(31);
	sub_wire2(193, 32)    <= sub_wire64(32);
	sub_wire2(193, 33)    <= sub_wire64(33);
	sub_wire2(193, 34)    <= sub_wire64(34);
	sub_wire2(193, 35)    <= sub_wire64(35);
	sub_wire2(193, 36)    <= sub_wire64(36);
	sub_wire2(193, 37)    <= sub_wire64(37);
	sub_wire2(193, 38)    <= sub_wire64(38);
	sub_wire2(193, 39)    <= sub_wire64(39);
	sub_wire2(192, 0)    <= sub_wire65(0);
	sub_wire2(192, 1)    <= sub_wire65(1);
	sub_wire2(192, 2)    <= sub_wire65(2);
	sub_wire2(192, 3)    <= sub_wire65(3);
	sub_wire2(192, 4)    <= sub_wire65(4);
	sub_wire2(192, 5)    <= sub_wire65(5);
	sub_wire2(192, 6)    <= sub_wire65(6);
	sub_wire2(192, 7)    <= sub_wire65(7);
	sub_wire2(192, 8)    <= sub_wire65(8);
	sub_wire2(192, 9)    <= sub_wire65(9);
	sub_wire2(192, 10)    <= sub_wire65(10);
	sub_wire2(192, 11)    <= sub_wire65(11);
	sub_wire2(192, 12)    <= sub_wire65(12);
	sub_wire2(192, 13)    <= sub_wire65(13);
	sub_wire2(192, 14)    <= sub_wire65(14);
	sub_wire2(192, 15)    <= sub_wire65(15);
	sub_wire2(192, 16)    <= sub_wire65(16);
	sub_wire2(192, 17)    <= sub_wire65(17);
	sub_wire2(192, 18)    <= sub_wire65(18);
	sub_wire2(192, 19)    <= sub_wire65(19);
	sub_wire2(192, 20)    <= sub_wire65(20);
	sub_wire2(192, 21)    <= sub_wire65(21);
	sub_wire2(192, 22)    <= sub_wire65(22);
	sub_wire2(192, 23)    <= sub_wire65(23);
	sub_wire2(192, 24)    <= sub_wire65(24);
	sub_wire2(192, 25)    <= sub_wire65(25);
	sub_wire2(192, 26)    <= sub_wire65(26);
	sub_wire2(192, 27)    <= sub_wire65(27);
	sub_wire2(192, 28)    <= sub_wire65(28);
	sub_wire2(192, 29)    <= sub_wire65(29);
	sub_wire2(192, 30)    <= sub_wire65(30);
	sub_wire2(192, 31)    <= sub_wire65(31);
	sub_wire2(192, 32)    <= sub_wire65(32);
	sub_wire2(192, 33)    <= sub_wire65(33);
	sub_wire2(192, 34)    <= sub_wire65(34);
	sub_wire2(192, 35)    <= sub_wire65(35);
	sub_wire2(192, 36)    <= sub_wire65(36);
	sub_wire2(192, 37)    <= sub_wire65(37);
	sub_wire2(192, 38)    <= sub_wire65(38);
	sub_wire2(192, 39)    <= sub_wire65(39);
	sub_wire2(191, 0)    <= sub_wire66(0);
	sub_wire2(191, 1)    <= sub_wire66(1);
	sub_wire2(191, 2)    <= sub_wire66(2);
	sub_wire2(191, 3)    <= sub_wire66(3);
	sub_wire2(191, 4)    <= sub_wire66(4);
	sub_wire2(191, 5)    <= sub_wire66(5);
	sub_wire2(191, 6)    <= sub_wire66(6);
	sub_wire2(191, 7)    <= sub_wire66(7);
	sub_wire2(191, 8)    <= sub_wire66(8);
	sub_wire2(191, 9)    <= sub_wire66(9);
	sub_wire2(191, 10)    <= sub_wire66(10);
	sub_wire2(191, 11)    <= sub_wire66(11);
	sub_wire2(191, 12)    <= sub_wire66(12);
	sub_wire2(191, 13)    <= sub_wire66(13);
	sub_wire2(191, 14)    <= sub_wire66(14);
	sub_wire2(191, 15)    <= sub_wire66(15);
	sub_wire2(191, 16)    <= sub_wire66(16);
	sub_wire2(191, 17)    <= sub_wire66(17);
	sub_wire2(191, 18)    <= sub_wire66(18);
	sub_wire2(191, 19)    <= sub_wire66(19);
	sub_wire2(191, 20)    <= sub_wire66(20);
	sub_wire2(191, 21)    <= sub_wire66(21);
	sub_wire2(191, 22)    <= sub_wire66(22);
	sub_wire2(191, 23)    <= sub_wire66(23);
	sub_wire2(191, 24)    <= sub_wire66(24);
	sub_wire2(191, 25)    <= sub_wire66(25);
	sub_wire2(191, 26)    <= sub_wire66(26);
	sub_wire2(191, 27)    <= sub_wire66(27);
	sub_wire2(191, 28)    <= sub_wire66(28);
	sub_wire2(191, 29)    <= sub_wire66(29);
	sub_wire2(191, 30)    <= sub_wire66(30);
	sub_wire2(191, 31)    <= sub_wire66(31);
	sub_wire2(191, 32)    <= sub_wire66(32);
	sub_wire2(191, 33)    <= sub_wire66(33);
	sub_wire2(191, 34)    <= sub_wire66(34);
	sub_wire2(191, 35)    <= sub_wire66(35);
	sub_wire2(191, 36)    <= sub_wire66(36);
	sub_wire2(191, 37)    <= sub_wire66(37);
	sub_wire2(191, 38)    <= sub_wire66(38);
	sub_wire2(191, 39)    <= sub_wire66(39);
	sub_wire2(190, 0)    <= sub_wire67(0);
	sub_wire2(190, 1)    <= sub_wire67(1);
	sub_wire2(190, 2)    <= sub_wire67(2);
	sub_wire2(190, 3)    <= sub_wire67(3);
	sub_wire2(190, 4)    <= sub_wire67(4);
	sub_wire2(190, 5)    <= sub_wire67(5);
	sub_wire2(190, 6)    <= sub_wire67(6);
	sub_wire2(190, 7)    <= sub_wire67(7);
	sub_wire2(190, 8)    <= sub_wire67(8);
	sub_wire2(190, 9)    <= sub_wire67(9);
	sub_wire2(190, 10)    <= sub_wire67(10);
	sub_wire2(190, 11)    <= sub_wire67(11);
	sub_wire2(190, 12)    <= sub_wire67(12);
	sub_wire2(190, 13)    <= sub_wire67(13);
	sub_wire2(190, 14)    <= sub_wire67(14);
	sub_wire2(190, 15)    <= sub_wire67(15);
	sub_wire2(190, 16)    <= sub_wire67(16);
	sub_wire2(190, 17)    <= sub_wire67(17);
	sub_wire2(190, 18)    <= sub_wire67(18);
	sub_wire2(190, 19)    <= sub_wire67(19);
	sub_wire2(190, 20)    <= sub_wire67(20);
	sub_wire2(190, 21)    <= sub_wire67(21);
	sub_wire2(190, 22)    <= sub_wire67(22);
	sub_wire2(190, 23)    <= sub_wire67(23);
	sub_wire2(190, 24)    <= sub_wire67(24);
	sub_wire2(190, 25)    <= sub_wire67(25);
	sub_wire2(190, 26)    <= sub_wire67(26);
	sub_wire2(190, 27)    <= sub_wire67(27);
	sub_wire2(190, 28)    <= sub_wire67(28);
	sub_wire2(190, 29)    <= sub_wire67(29);
	sub_wire2(190, 30)    <= sub_wire67(30);
	sub_wire2(190, 31)    <= sub_wire67(31);
	sub_wire2(190, 32)    <= sub_wire67(32);
	sub_wire2(190, 33)    <= sub_wire67(33);
	sub_wire2(190, 34)    <= sub_wire67(34);
	sub_wire2(190, 35)    <= sub_wire67(35);
	sub_wire2(190, 36)    <= sub_wire67(36);
	sub_wire2(190, 37)    <= sub_wire67(37);
	sub_wire2(190, 38)    <= sub_wire67(38);
	sub_wire2(190, 39)    <= sub_wire67(39);
	sub_wire2(189, 0)    <= sub_wire68(0);
	sub_wire2(189, 1)    <= sub_wire68(1);
	sub_wire2(189, 2)    <= sub_wire68(2);
	sub_wire2(189, 3)    <= sub_wire68(3);
	sub_wire2(189, 4)    <= sub_wire68(4);
	sub_wire2(189, 5)    <= sub_wire68(5);
	sub_wire2(189, 6)    <= sub_wire68(6);
	sub_wire2(189, 7)    <= sub_wire68(7);
	sub_wire2(189, 8)    <= sub_wire68(8);
	sub_wire2(189, 9)    <= sub_wire68(9);
	sub_wire2(189, 10)    <= sub_wire68(10);
	sub_wire2(189, 11)    <= sub_wire68(11);
	sub_wire2(189, 12)    <= sub_wire68(12);
	sub_wire2(189, 13)    <= sub_wire68(13);
	sub_wire2(189, 14)    <= sub_wire68(14);
	sub_wire2(189, 15)    <= sub_wire68(15);
	sub_wire2(189, 16)    <= sub_wire68(16);
	sub_wire2(189, 17)    <= sub_wire68(17);
	sub_wire2(189, 18)    <= sub_wire68(18);
	sub_wire2(189, 19)    <= sub_wire68(19);
	sub_wire2(189, 20)    <= sub_wire68(20);
	sub_wire2(189, 21)    <= sub_wire68(21);
	sub_wire2(189, 22)    <= sub_wire68(22);
	sub_wire2(189, 23)    <= sub_wire68(23);
	sub_wire2(189, 24)    <= sub_wire68(24);
	sub_wire2(189, 25)    <= sub_wire68(25);
	sub_wire2(189, 26)    <= sub_wire68(26);
	sub_wire2(189, 27)    <= sub_wire68(27);
	sub_wire2(189, 28)    <= sub_wire68(28);
	sub_wire2(189, 29)    <= sub_wire68(29);
	sub_wire2(189, 30)    <= sub_wire68(30);
	sub_wire2(189, 31)    <= sub_wire68(31);
	sub_wire2(189, 32)    <= sub_wire68(32);
	sub_wire2(189, 33)    <= sub_wire68(33);
	sub_wire2(189, 34)    <= sub_wire68(34);
	sub_wire2(189, 35)    <= sub_wire68(35);
	sub_wire2(189, 36)    <= sub_wire68(36);
	sub_wire2(189, 37)    <= sub_wire68(37);
	sub_wire2(189, 38)    <= sub_wire68(38);
	sub_wire2(189, 39)    <= sub_wire68(39);
	sub_wire2(188, 0)    <= sub_wire69(0);
	sub_wire2(188, 1)    <= sub_wire69(1);
	sub_wire2(188, 2)    <= sub_wire69(2);
	sub_wire2(188, 3)    <= sub_wire69(3);
	sub_wire2(188, 4)    <= sub_wire69(4);
	sub_wire2(188, 5)    <= sub_wire69(5);
	sub_wire2(188, 6)    <= sub_wire69(6);
	sub_wire2(188, 7)    <= sub_wire69(7);
	sub_wire2(188, 8)    <= sub_wire69(8);
	sub_wire2(188, 9)    <= sub_wire69(9);
	sub_wire2(188, 10)    <= sub_wire69(10);
	sub_wire2(188, 11)    <= sub_wire69(11);
	sub_wire2(188, 12)    <= sub_wire69(12);
	sub_wire2(188, 13)    <= sub_wire69(13);
	sub_wire2(188, 14)    <= sub_wire69(14);
	sub_wire2(188, 15)    <= sub_wire69(15);
	sub_wire2(188, 16)    <= sub_wire69(16);
	sub_wire2(188, 17)    <= sub_wire69(17);
	sub_wire2(188, 18)    <= sub_wire69(18);
	sub_wire2(188, 19)    <= sub_wire69(19);
	sub_wire2(188, 20)    <= sub_wire69(20);
	sub_wire2(188, 21)    <= sub_wire69(21);
	sub_wire2(188, 22)    <= sub_wire69(22);
	sub_wire2(188, 23)    <= sub_wire69(23);
	sub_wire2(188, 24)    <= sub_wire69(24);
	sub_wire2(188, 25)    <= sub_wire69(25);
	sub_wire2(188, 26)    <= sub_wire69(26);
	sub_wire2(188, 27)    <= sub_wire69(27);
	sub_wire2(188, 28)    <= sub_wire69(28);
	sub_wire2(188, 29)    <= sub_wire69(29);
	sub_wire2(188, 30)    <= sub_wire69(30);
	sub_wire2(188, 31)    <= sub_wire69(31);
	sub_wire2(188, 32)    <= sub_wire69(32);
	sub_wire2(188, 33)    <= sub_wire69(33);
	sub_wire2(188, 34)    <= sub_wire69(34);
	sub_wire2(188, 35)    <= sub_wire69(35);
	sub_wire2(188, 36)    <= sub_wire69(36);
	sub_wire2(188, 37)    <= sub_wire69(37);
	sub_wire2(188, 38)    <= sub_wire69(38);
	sub_wire2(188, 39)    <= sub_wire69(39);
	sub_wire2(187, 0)    <= sub_wire70(0);
	sub_wire2(187, 1)    <= sub_wire70(1);
	sub_wire2(187, 2)    <= sub_wire70(2);
	sub_wire2(187, 3)    <= sub_wire70(3);
	sub_wire2(187, 4)    <= sub_wire70(4);
	sub_wire2(187, 5)    <= sub_wire70(5);
	sub_wire2(187, 6)    <= sub_wire70(6);
	sub_wire2(187, 7)    <= sub_wire70(7);
	sub_wire2(187, 8)    <= sub_wire70(8);
	sub_wire2(187, 9)    <= sub_wire70(9);
	sub_wire2(187, 10)    <= sub_wire70(10);
	sub_wire2(187, 11)    <= sub_wire70(11);
	sub_wire2(187, 12)    <= sub_wire70(12);
	sub_wire2(187, 13)    <= sub_wire70(13);
	sub_wire2(187, 14)    <= sub_wire70(14);
	sub_wire2(187, 15)    <= sub_wire70(15);
	sub_wire2(187, 16)    <= sub_wire70(16);
	sub_wire2(187, 17)    <= sub_wire70(17);
	sub_wire2(187, 18)    <= sub_wire70(18);
	sub_wire2(187, 19)    <= sub_wire70(19);
	sub_wire2(187, 20)    <= sub_wire70(20);
	sub_wire2(187, 21)    <= sub_wire70(21);
	sub_wire2(187, 22)    <= sub_wire70(22);
	sub_wire2(187, 23)    <= sub_wire70(23);
	sub_wire2(187, 24)    <= sub_wire70(24);
	sub_wire2(187, 25)    <= sub_wire70(25);
	sub_wire2(187, 26)    <= sub_wire70(26);
	sub_wire2(187, 27)    <= sub_wire70(27);
	sub_wire2(187, 28)    <= sub_wire70(28);
	sub_wire2(187, 29)    <= sub_wire70(29);
	sub_wire2(187, 30)    <= sub_wire70(30);
	sub_wire2(187, 31)    <= sub_wire70(31);
	sub_wire2(187, 32)    <= sub_wire70(32);
	sub_wire2(187, 33)    <= sub_wire70(33);
	sub_wire2(187, 34)    <= sub_wire70(34);
	sub_wire2(187, 35)    <= sub_wire70(35);
	sub_wire2(187, 36)    <= sub_wire70(36);
	sub_wire2(187, 37)    <= sub_wire70(37);
	sub_wire2(187, 38)    <= sub_wire70(38);
	sub_wire2(187, 39)    <= sub_wire70(39);
	sub_wire2(186, 0)    <= sub_wire71(0);
	sub_wire2(186, 1)    <= sub_wire71(1);
	sub_wire2(186, 2)    <= sub_wire71(2);
	sub_wire2(186, 3)    <= sub_wire71(3);
	sub_wire2(186, 4)    <= sub_wire71(4);
	sub_wire2(186, 5)    <= sub_wire71(5);
	sub_wire2(186, 6)    <= sub_wire71(6);
	sub_wire2(186, 7)    <= sub_wire71(7);
	sub_wire2(186, 8)    <= sub_wire71(8);
	sub_wire2(186, 9)    <= sub_wire71(9);
	sub_wire2(186, 10)    <= sub_wire71(10);
	sub_wire2(186, 11)    <= sub_wire71(11);
	sub_wire2(186, 12)    <= sub_wire71(12);
	sub_wire2(186, 13)    <= sub_wire71(13);
	sub_wire2(186, 14)    <= sub_wire71(14);
	sub_wire2(186, 15)    <= sub_wire71(15);
	sub_wire2(186, 16)    <= sub_wire71(16);
	sub_wire2(186, 17)    <= sub_wire71(17);
	sub_wire2(186, 18)    <= sub_wire71(18);
	sub_wire2(186, 19)    <= sub_wire71(19);
	sub_wire2(186, 20)    <= sub_wire71(20);
	sub_wire2(186, 21)    <= sub_wire71(21);
	sub_wire2(186, 22)    <= sub_wire71(22);
	sub_wire2(186, 23)    <= sub_wire71(23);
	sub_wire2(186, 24)    <= sub_wire71(24);
	sub_wire2(186, 25)    <= sub_wire71(25);
	sub_wire2(186, 26)    <= sub_wire71(26);
	sub_wire2(186, 27)    <= sub_wire71(27);
	sub_wire2(186, 28)    <= sub_wire71(28);
	sub_wire2(186, 29)    <= sub_wire71(29);
	sub_wire2(186, 30)    <= sub_wire71(30);
	sub_wire2(186, 31)    <= sub_wire71(31);
	sub_wire2(186, 32)    <= sub_wire71(32);
	sub_wire2(186, 33)    <= sub_wire71(33);
	sub_wire2(186, 34)    <= sub_wire71(34);
	sub_wire2(186, 35)    <= sub_wire71(35);
	sub_wire2(186, 36)    <= sub_wire71(36);
	sub_wire2(186, 37)    <= sub_wire71(37);
	sub_wire2(186, 38)    <= sub_wire71(38);
	sub_wire2(186, 39)    <= sub_wire71(39);
	sub_wire2(185, 0)    <= sub_wire72(0);
	sub_wire2(185, 1)    <= sub_wire72(1);
	sub_wire2(185, 2)    <= sub_wire72(2);
	sub_wire2(185, 3)    <= sub_wire72(3);
	sub_wire2(185, 4)    <= sub_wire72(4);
	sub_wire2(185, 5)    <= sub_wire72(5);
	sub_wire2(185, 6)    <= sub_wire72(6);
	sub_wire2(185, 7)    <= sub_wire72(7);
	sub_wire2(185, 8)    <= sub_wire72(8);
	sub_wire2(185, 9)    <= sub_wire72(9);
	sub_wire2(185, 10)    <= sub_wire72(10);
	sub_wire2(185, 11)    <= sub_wire72(11);
	sub_wire2(185, 12)    <= sub_wire72(12);
	sub_wire2(185, 13)    <= sub_wire72(13);
	sub_wire2(185, 14)    <= sub_wire72(14);
	sub_wire2(185, 15)    <= sub_wire72(15);
	sub_wire2(185, 16)    <= sub_wire72(16);
	sub_wire2(185, 17)    <= sub_wire72(17);
	sub_wire2(185, 18)    <= sub_wire72(18);
	sub_wire2(185, 19)    <= sub_wire72(19);
	sub_wire2(185, 20)    <= sub_wire72(20);
	sub_wire2(185, 21)    <= sub_wire72(21);
	sub_wire2(185, 22)    <= sub_wire72(22);
	sub_wire2(185, 23)    <= sub_wire72(23);
	sub_wire2(185, 24)    <= sub_wire72(24);
	sub_wire2(185, 25)    <= sub_wire72(25);
	sub_wire2(185, 26)    <= sub_wire72(26);
	sub_wire2(185, 27)    <= sub_wire72(27);
	sub_wire2(185, 28)    <= sub_wire72(28);
	sub_wire2(185, 29)    <= sub_wire72(29);
	sub_wire2(185, 30)    <= sub_wire72(30);
	sub_wire2(185, 31)    <= sub_wire72(31);
	sub_wire2(185, 32)    <= sub_wire72(32);
	sub_wire2(185, 33)    <= sub_wire72(33);
	sub_wire2(185, 34)    <= sub_wire72(34);
	sub_wire2(185, 35)    <= sub_wire72(35);
	sub_wire2(185, 36)    <= sub_wire72(36);
	sub_wire2(185, 37)    <= sub_wire72(37);
	sub_wire2(185, 38)    <= sub_wire72(38);
	sub_wire2(185, 39)    <= sub_wire72(39);
	sub_wire2(184, 0)    <= sub_wire73(0);
	sub_wire2(184, 1)    <= sub_wire73(1);
	sub_wire2(184, 2)    <= sub_wire73(2);
	sub_wire2(184, 3)    <= sub_wire73(3);
	sub_wire2(184, 4)    <= sub_wire73(4);
	sub_wire2(184, 5)    <= sub_wire73(5);
	sub_wire2(184, 6)    <= sub_wire73(6);
	sub_wire2(184, 7)    <= sub_wire73(7);
	sub_wire2(184, 8)    <= sub_wire73(8);
	sub_wire2(184, 9)    <= sub_wire73(9);
	sub_wire2(184, 10)    <= sub_wire73(10);
	sub_wire2(184, 11)    <= sub_wire73(11);
	sub_wire2(184, 12)    <= sub_wire73(12);
	sub_wire2(184, 13)    <= sub_wire73(13);
	sub_wire2(184, 14)    <= sub_wire73(14);
	sub_wire2(184, 15)    <= sub_wire73(15);
	sub_wire2(184, 16)    <= sub_wire73(16);
	sub_wire2(184, 17)    <= sub_wire73(17);
	sub_wire2(184, 18)    <= sub_wire73(18);
	sub_wire2(184, 19)    <= sub_wire73(19);
	sub_wire2(184, 20)    <= sub_wire73(20);
	sub_wire2(184, 21)    <= sub_wire73(21);
	sub_wire2(184, 22)    <= sub_wire73(22);
	sub_wire2(184, 23)    <= sub_wire73(23);
	sub_wire2(184, 24)    <= sub_wire73(24);
	sub_wire2(184, 25)    <= sub_wire73(25);
	sub_wire2(184, 26)    <= sub_wire73(26);
	sub_wire2(184, 27)    <= sub_wire73(27);
	sub_wire2(184, 28)    <= sub_wire73(28);
	sub_wire2(184, 29)    <= sub_wire73(29);
	sub_wire2(184, 30)    <= sub_wire73(30);
	sub_wire2(184, 31)    <= sub_wire73(31);
	sub_wire2(184, 32)    <= sub_wire73(32);
	sub_wire2(184, 33)    <= sub_wire73(33);
	sub_wire2(184, 34)    <= sub_wire73(34);
	sub_wire2(184, 35)    <= sub_wire73(35);
	sub_wire2(184, 36)    <= sub_wire73(36);
	sub_wire2(184, 37)    <= sub_wire73(37);
	sub_wire2(184, 38)    <= sub_wire73(38);
	sub_wire2(184, 39)    <= sub_wire73(39);
	sub_wire2(183, 0)    <= sub_wire74(0);
	sub_wire2(183, 1)    <= sub_wire74(1);
	sub_wire2(183, 2)    <= sub_wire74(2);
	sub_wire2(183, 3)    <= sub_wire74(3);
	sub_wire2(183, 4)    <= sub_wire74(4);
	sub_wire2(183, 5)    <= sub_wire74(5);
	sub_wire2(183, 6)    <= sub_wire74(6);
	sub_wire2(183, 7)    <= sub_wire74(7);
	sub_wire2(183, 8)    <= sub_wire74(8);
	sub_wire2(183, 9)    <= sub_wire74(9);
	sub_wire2(183, 10)    <= sub_wire74(10);
	sub_wire2(183, 11)    <= sub_wire74(11);
	sub_wire2(183, 12)    <= sub_wire74(12);
	sub_wire2(183, 13)    <= sub_wire74(13);
	sub_wire2(183, 14)    <= sub_wire74(14);
	sub_wire2(183, 15)    <= sub_wire74(15);
	sub_wire2(183, 16)    <= sub_wire74(16);
	sub_wire2(183, 17)    <= sub_wire74(17);
	sub_wire2(183, 18)    <= sub_wire74(18);
	sub_wire2(183, 19)    <= sub_wire74(19);
	sub_wire2(183, 20)    <= sub_wire74(20);
	sub_wire2(183, 21)    <= sub_wire74(21);
	sub_wire2(183, 22)    <= sub_wire74(22);
	sub_wire2(183, 23)    <= sub_wire74(23);
	sub_wire2(183, 24)    <= sub_wire74(24);
	sub_wire2(183, 25)    <= sub_wire74(25);
	sub_wire2(183, 26)    <= sub_wire74(26);
	sub_wire2(183, 27)    <= sub_wire74(27);
	sub_wire2(183, 28)    <= sub_wire74(28);
	sub_wire2(183, 29)    <= sub_wire74(29);
	sub_wire2(183, 30)    <= sub_wire74(30);
	sub_wire2(183, 31)    <= sub_wire74(31);
	sub_wire2(183, 32)    <= sub_wire74(32);
	sub_wire2(183, 33)    <= sub_wire74(33);
	sub_wire2(183, 34)    <= sub_wire74(34);
	sub_wire2(183, 35)    <= sub_wire74(35);
	sub_wire2(183, 36)    <= sub_wire74(36);
	sub_wire2(183, 37)    <= sub_wire74(37);
	sub_wire2(183, 38)    <= sub_wire74(38);
	sub_wire2(183, 39)    <= sub_wire74(39);
	sub_wire2(182, 0)    <= sub_wire75(0);
	sub_wire2(182, 1)    <= sub_wire75(1);
	sub_wire2(182, 2)    <= sub_wire75(2);
	sub_wire2(182, 3)    <= sub_wire75(3);
	sub_wire2(182, 4)    <= sub_wire75(4);
	sub_wire2(182, 5)    <= sub_wire75(5);
	sub_wire2(182, 6)    <= sub_wire75(6);
	sub_wire2(182, 7)    <= sub_wire75(7);
	sub_wire2(182, 8)    <= sub_wire75(8);
	sub_wire2(182, 9)    <= sub_wire75(9);
	sub_wire2(182, 10)    <= sub_wire75(10);
	sub_wire2(182, 11)    <= sub_wire75(11);
	sub_wire2(182, 12)    <= sub_wire75(12);
	sub_wire2(182, 13)    <= sub_wire75(13);
	sub_wire2(182, 14)    <= sub_wire75(14);
	sub_wire2(182, 15)    <= sub_wire75(15);
	sub_wire2(182, 16)    <= sub_wire75(16);
	sub_wire2(182, 17)    <= sub_wire75(17);
	sub_wire2(182, 18)    <= sub_wire75(18);
	sub_wire2(182, 19)    <= sub_wire75(19);
	sub_wire2(182, 20)    <= sub_wire75(20);
	sub_wire2(182, 21)    <= sub_wire75(21);
	sub_wire2(182, 22)    <= sub_wire75(22);
	sub_wire2(182, 23)    <= sub_wire75(23);
	sub_wire2(182, 24)    <= sub_wire75(24);
	sub_wire2(182, 25)    <= sub_wire75(25);
	sub_wire2(182, 26)    <= sub_wire75(26);
	sub_wire2(182, 27)    <= sub_wire75(27);
	sub_wire2(182, 28)    <= sub_wire75(28);
	sub_wire2(182, 29)    <= sub_wire75(29);
	sub_wire2(182, 30)    <= sub_wire75(30);
	sub_wire2(182, 31)    <= sub_wire75(31);
	sub_wire2(182, 32)    <= sub_wire75(32);
	sub_wire2(182, 33)    <= sub_wire75(33);
	sub_wire2(182, 34)    <= sub_wire75(34);
	sub_wire2(182, 35)    <= sub_wire75(35);
	sub_wire2(182, 36)    <= sub_wire75(36);
	sub_wire2(182, 37)    <= sub_wire75(37);
	sub_wire2(182, 38)    <= sub_wire75(38);
	sub_wire2(182, 39)    <= sub_wire75(39);
	sub_wire2(181, 0)    <= sub_wire76(0);
	sub_wire2(181, 1)    <= sub_wire76(1);
	sub_wire2(181, 2)    <= sub_wire76(2);
	sub_wire2(181, 3)    <= sub_wire76(3);
	sub_wire2(181, 4)    <= sub_wire76(4);
	sub_wire2(181, 5)    <= sub_wire76(5);
	sub_wire2(181, 6)    <= sub_wire76(6);
	sub_wire2(181, 7)    <= sub_wire76(7);
	sub_wire2(181, 8)    <= sub_wire76(8);
	sub_wire2(181, 9)    <= sub_wire76(9);
	sub_wire2(181, 10)    <= sub_wire76(10);
	sub_wire2(181, 11)    <= sub_wire76(11);
	sub_wire2(181, 12)    <= sub_wire76(12);
	sub_wire2(181, 13)    <= sub_wire76(13);
	sub_wire2(181, 14)    <= sub_wire76(14);
	sub_wire2(181, 15)    <= sub_wire76(15);
	sub_wire2(181, 16)    <= sub_wire76(16);
	sub_wire2(181, 17)    <= sub_wire76(17);
	sub_wire2(181, 18)    <= sub_wire76(18);
	sub_wire2(181, 19)    <= sub_wire76(19);
	sub_wire2(181, 20)    <= sub_wire76(20);
	sub_wire2(181, 21)    <= sub_wire76(21);
	sub_wire2(181, 22)    <= sub_wire76(22);
	sub_wire2(181, 23)    <= sub_wire76(23);
	sub_wire2(181, 24)    <= sub_wire76(24);
	sub_wire2(181, 25)    <= sub_wire76(25);
	sub_wire2(181, 26)    <= sub_wire76(26);
	sub_wire2(181, 27)    <= sub_wire76(27);
	sub_wire2(181, 28)    <= sub_wire76(28);
	sub_wire2(181, 29)    <= sub_wire76(29);
	sub_wire2(181, 30)    <= sub_wire76(30);
	sub_wire2(181, 31)    <= sub_wire76(31);
	sub_wire2(181, 32)    <= sub_wire76(32);
	sub_wire2(181, 33)    <= sub_wire76(33);
	sub_wire2(181, 34)    <= sub_wire76(34);
	sub_wire2(181, 35)    <= sub_wire76(35);
	sub_wire2(181, 36)    <= sub_wire76(36);
	sub_wire2(181, 37)    <= sub_wire76(37);
	sub_wire2(181, 38)    <= sub_wire76(38);
	sub_wire2(181, 39)    <= sub_wire76(39);
	sub_wire2(180, 0)    <= sub_wire77(0);
	sub_wire2(180, 1)    <= sub_wire77(1);
	sub_wire2(180, 2)    <= sub_wire77(2);
	sub_wire2(180, 3)    <= sub_wire77(3);
	sub_wire2(180, 4)    <= sub_wire77(4);
	sub_wire2(180, 5)    <= sub_wire77(5);
	sub_wire2(180, 6)    <= sub_wire77(6);
	sub_wire2(180, 7)    <= sub_wire77(7);
	sub_wire2(180, 8)    <= sub_wire77(8);
	sub_wire2(180, 9)    <= sub_wire77(9);
	sub_wire2(180, 10)    <= sub_wire77(10);
	sub_wire2(180, 11)    <= sub_wire77(11);
	sub_wire2(180, 12)    <= sub_wire77(12);
	sub_wire2(180, 13)    <= sub_wire77(13);
	sub_wire2(180, 14)    <= sub_wire77(14);
	sub_wire2(180, 15)    <= sub_wire77(15);
	sub_wire2(180, 16)    <= sub_wire77(16);
	sub_wire2(180, 17)    <= sub_wire77(17);
	sub_wire2(180, 18)    <= sub_wire77(18);
	sub_wire2(180, 19)    <= sub_wire77(19);
	sub_wire2(180, 20)    <= sub_wire77(20);
	sub_wire2(180, 21)    <= sub_wire77(21);
	sub_wire2(180, 22)    <= sub_wire77(22);
	sub_wire2(180, 23)    <= sub_wire77(23);
	sub_wire2(180, 24)    <= sub_wire77(24);
	sub_wire2(180, 25)    <= sub_wire77(25);
	sub_wire2(180, 26)    <= sub_wire77(26);
	sub_wire2(180, 27)    <= sub_wire77(27);
	sub_wire2(180, 28)    <= sub_wire77(28);
	sub_wire2(180, 29)    <= sub_wire77(29);
	sub_wire2(180, 30)    <= sub_wire77(30);
	sub_wire2(180, 31)    <= sub_wire77(31);
	sub_wire2(180, 32)    <= sub_wire77(32);
	sub_wire2(180, 33)    <= sub_wire77(33);
	sub_wire2(180, 34)    <= sub_wire77(34);
	sub_wire2(180, 35)    <= sub_wire77(35);
	sub_wire2(180, 36)    <= sub_wire77(36);
	sub_wire2(180, 37)    <= sub_wire77(37);
	sub_wire2(180, 38)    <= sub_wire77(38);
	sub_wire2(180, 39)    <= sub_wire77(39);
	sub_wire2(179, 0)    <= sub_wire78(0);
	sub_wire2(179, 1)    <= sub_wire78(1);
	sub_wire2(179, 2)    <= sub_wire78(2);
	sub_wire2(179, 3)    <= sub_wire78(3);
	sub_wire2(179, 4)    <= sub_wire78(4);
	sub_wire2(179, 5)    <= sub_wire78(5);
	sub_wire2(179, 6)    <= sub_wire78(6);
	sub_wire2(179, 7)    <= sub_wire78(7);
	sub_wire2(179, 8)    <= sub_wire78(8);
	sub_wire2(179, 9)    <= sub_wire78(9);
	sub_wire2(179, 10)    <= sub_wire78(10);
	sub_wire2(179, 11)    <= sub_wire78(11);
	sub_wire2(179, 12)    <= sub_wire78(12);
	sub_wire2(179, 13)    <= sub_wire78(13);
	sub_wire2(179, 14)    <= sub_wire78(14);
	sub_wire2(179, 15)    <= sub_wire78(15);
	sub_wire2(179, 16)    <= sub_wire78(16);
	sub_wire2(179, 17)    <= sub_wire78(17);
	sub_wire2(179, 18)    <= sub_wire78(18);
	sub_wire2(179, 19)    <= sub_wire78(19);
	sub_wire2(179, 20)    <= sub_wire78(20);
	sub_wire2(179, 21)    <= sub_wire78(21);
	sub_wire2(179, 22)    <= sub_wire78(22);
	sub_wire2(179, 23)    <= sub_wire78(23);
	sub_wire2(179, 24)    <= sub_wire78(24);
	sub_wire2(179, 25)    <= sub_wire78(25);
	sub_wire2(179, 26)    <= sub_wire78(26);
	sub_wire2(179, 27)    <= sub_wire78(27);
	sub_wire2(179, 28)    <= sub_wire78(28);
	sub_wire2(179, 29)    <= sub_wire78(29);
	sub_wire2(179, 30)    <= sub_wire78(30);
	sub_wire2(179, 31)    <= sub_wire78(31);
	sub_wire2(179, 32)    <= sub_wire78(32);
	sub_wire2(179, 33)    <= sub_wire78(33);
	sub_wire2(179, 34)    <= sub_wire78(34);
	sub_wire2(179, 35)    <= sub_wire78(35);
	sub_wire2(179, 36)    <= sub_wire78(36);
	sub_wire2(179, 37)    <= sub_wire78(37);
	sub_wire2(179, 38)    <= sub_wire78(38);
	sub_wire2(179, 39)    <= sub_wire78(39);
	sub_wire2(178, 0)    <= sub_wire79(0);
	sub_wire2(178, 1)    <= sub_wire79(1);
	sub_wire2(178, 2)    <= sub_wire79(2);
	sub_wire2(178, 3)    <= sub_wire79(3);
	sub_wire2(178, 4)    <= sub_wire79(4);
	sub_wire2(178, 5)    <= sub_wire79(5);
	sub_wire2(178, 6)    <= sub_wire79(6);
	sub_wire2(178, 7)    <= sub_wire79(7);
	sub_wire2(178, 8)    <= sub_wire79(8);
	sub_wire2(178, 9)    <= sub_wire79(9);
	sub_wire2(178, 10)    <= sub_wire79(10);
	sub_wire2(178, 11)    <= sub_wire79(11);
	sub_wire2(178, 12)    <= sub_wire79(12);
	sub_wire2(178, 13)    <= sub_wire79(13);
	sub_wire2(178, 14)    <= sub_wire79(14);
	sub_wire2(178, 15)    <= sub_wire79(15);
	sub_wire2(178, 16)    <= sub_wire79(16);
	sub_wire2(178, 17)    <= sub_wire79(17);
	sub_wire2(178, 18)    <= sub_wire79(18);
	sub_wire2(178, 19)    <= sub_wire79(19);
	sub_wire2(178, 20)    <= sub_wire79(20);
	sub_wire2(178, 21)    <= sub_wire79(21);
	sub_wire2(178, 22)    <= sub_wire79(22);
	sub_wire2(178, 23)    <= sub_wire79(23);
	sub_wire2(178, 24)    <= sub_wire79(24);
	sub_wire2(178, 25)    <= sub_wire79(25);
	sub_wire2(178, 26)    <= sub_wire79(26);
	sub_wire2(178, 27)    <= sub_wire79(27);
	sub_wire2(178, 28)    <= sub_wire79(28);
	sub_wire2(178, 29)    <= sub_wire79(29);
	sub_wire2(178, 30)    <= sub_wire79(30);
	sub_wire2(178, 31)    <= sub_wire79(31);
	sub_wire2(178, 32)    <= sub_wire79(32);
	sub_wire2(178, 33)    <= sub_wire79(33);
	sub_wire2(178, 34)    <= sub_wire79(34);
	sub_wire2(178, 35)    <= sub_wire79(35);
	sub_wire2(178, 36)    <= sub_wire79(36);
	sub_wire2(178, 37)    <= sub_wire79(37);
	sub_wire2(178, 38)    <= sub_wire79(38);
	sub_wire2(178, 39)    <= sub_wire79(39);
	sub_wire2(177, 0)    <= sub_wire80(0);
	sub_wire2(177, 1)    <= sub_wire80(1);
	sub_wire2(177, 2)    <= sub_wire80(2);
	sub_wire2(177, 3)    <= sub_wire80(3);
	sub_wire2(177, 4)    <= sub_wire80(4);
	sub_wire2(177, 5)    <= sub_wire80(5);
	sub_wire2(177, 6)    <= sub_wire80(6);
	sub_wire2(177, 7)    <= sub_wire80(7);
	sub_wire2(177, 8)    <= sub_wire80(8);
	sub_wire2(177, 9)    <= sub_wire80(9);
	sub_wire2(177, 10)    <= sub_wire80(10);
	sub_wire2(177, 11)    <= sub_wire80(11);
	sub_wire2(177, 12)    <= sub_wire80(12);
	sub_wire2(177, 13)    <= sub_wire80(13);
	sub_wire2(177, 14)    <= sub_wire80(14);
	sub_wire2(177, 15)    <= sub_wire80(15);
	sub_wire2(177, 16)    <= sub_wire80(16);
	sub_wire2(177, 17)    <= sub_wire80(17);
	sub_wire2(177, 18)    <= sub_wire80(18);
	sub_wire2(177, 19)    <= sub_wire80(19);
	sub_wire2(177, 20)    <= sub_wire80(20);
	sub_wire2(177, 21)    <= sub_wire80(21);
	sub_wire2(177, 22)    <= sub_wire80(22);
	sub_wire2(177, 23)    <= sub_wire80(23);
	sub_wire2(177, 24)    <= sub_wire80(24);
	sub_wire2(177, 25)    <= sub_wire80(25);
	sub_wire2(177, 26)    <= sub_wire80(26);
	sub_wire2(177, 27)    <= sub_wire80(27);
	sub_wire2(177, 28)    <= sub_wire80(28);
	sub_wire2(177, 29)    <= sub_wire80(29);
	sub_wire2(177, 30)    <= sub_wire80(30);
	sub_wire2(177, 31)    <= sub_wire80(31);
	sub_wire2(177, 32)    <= sub_wire80(32);
	sub_wire2(177, 33)    <= sub_wire80(33);
	sub_wire2(177, 34)    <= sub_wire80(34);
	sub_wire2(177, 35)    <= sub_wire80(35);
	sub_wire2(177, 36)    <= sub_wire80(36);
	sub_wire2(177, 37)    <= sub_wire80(37);
	sub_wire2(177, 38)    <= sub_wire80(38);
	sub_wire2(177, 39)    <= sub_wire80(39);
	sub_wire2(176, 0)    <= sub_wire81(0);
	sub_wire2(176, 1)    <= sub_wire81(1);
	sub_wire2(176, 2)    <= sub_wire81(2);
	sub_wire2(176, 3)    <= sub_wire81(3);
	sub_wire2(176, 4)    <= sub_wire81(4);
	sub_wire2(176, 5)    <= sub_wire81(5);
	sub_wire2(176, 6)    <= sub_wire81(6);
	sub_wire2(176, 7)    <= sub_wire81(7);
	sub_wire2(176, 8)    <= sub_wire81(8);
	sub_wire2(176, 9)    <= sub_wire81(9);
	sub_wire2(176, 10)    <= sub_wire81(10);
	sub_wire2(176, 11)    <= sub_wire81(11);
	sub_wire2(176, 12)    <= sub_wire81(12);
	sub_wire2(176, 13)    <= sub_wire81(13);
	sub_wire2(176, 14)    <= sub_wire81(14);
	sub_wire2(176, 15)    <= sub_wire81(15);
	sub_wire2(176, 16)    <= sub_wire81(16);
	sub_wire2(176, 17)    <= sub_wire81(17);
	sub_wire2(176, 18)    <= sub_wire81(18);
	sub_wire2(176, 19)    <= sub_wire81(19);
	sub_wire2(176, 20)    <= sub_wire81(20);
	sub_wire2(176, 21)    <= sub_wire81(21);
	sub_wire2(176, 22)    <= sub_wire81(22);
	sub_wire2(176, 23)    <= sub_wire81(23);
	sub_wire2(176, 24)    <= sub_wire81(24);
	sub_wire2(176, 25)    <= sub_wire81(25);
	sub_wire2(176, 26)    <= sub_wire81(26);
	sub_wire2(176, 27)    <= sub_wire81(27);
	sub_wire2(176, 28)    <= sub_wire81(28);
	sub_wire2(176, 29)    <= sub_wire81(29);
	sub_wire2(176, 30)    <= sub_wire81(30);
	sub_wire2(176, 31)    <= sub_wire81(31);
	sub_wire2(176, 32)    <= sub_wire81(32);
	sub_wire2(176, 33)    <= sub_wire81(33);
	sub_wire2(176, 34)    <= sub_wire81(34);
	sub_wire2(176, 35)    <= sub_wire81(35);
	sub_wire2(176, 36)    <= sub_wire81(36);
	sub_wire2(176, 37)    <= sub_wire81(37);
	sub_wire2(176, 38)    <= sub_wire81(38);
	sub_wire2(176, 39)    <= sub_wire81(39);
	sub_wire2(175, 0)    <= sub_wire82(0);
	sub_wire2(175, 1)    <= sub_wire82(1);
	sub_wire2(175, 2)    <= sub_wire82(2);
	sub_wire2(175, 3)    <= sub_wire82(3);
	sub_wire2(175, 4)    <= sub_wire82(4);
	sub_wire2(175, 5)    <= sub_wire82(5);
	sub_wire2(175, 6)    <= sub_wire82(6);
	sub_wire2(175, 7)    <= sub_wire82(7);
	sub_wire2(175, 8)    <= sub_wire82(8);
	sub_wire2(175, 9)    <= sub_wire82(9);
	sub_wire2(175, 10)    <= sub_wire82(10);
	sub_wire2(175, 11)    <= sub_wire82(11);
	sub_wire2(175, 12)    <= sub_wire82(12);
	sub_wire2(175, 13)    <= sub_wire82(13);
	sub_wire2(175, 14)    <= sub_wire82(14);
	sub_wire2(175, 15)    <= sub_wire82(15);
	sub_wire2(175, 16)    <= sub_wire82(16);
	sub_wire2(175, 17)    <= sub_wire82(17);
	sub_wire2(175, 18)    <= sub_wire82(18);
	sub_wire2(175, 19)    <= sub_wire82(19);
	sub_wire2(175, 20)    <= sub_wire82(20);
	sub_wire2(175, 21)    <= sub_wire82(21);
	sub_wire2(175, 22)    <= sub_wire82(22);
	sub_wire2(175, 23)    <= sub_wire82(23);
	sub_wire2(175, 24)    <= sub_wire82(24);
	sub_wire2(175, 25)    <= sub_wire82(25);
	sub_wire2(175, 26)    <= sub_wire82(26);
	sub_wire2(175, 27)    <= sub_wire82(27);
	sub_wire2(175, 28)    <= sub_wire82(28);
	sub_wire2(175, 29)    <= sub_wire82(29);
	sub_wire2(175, 30)    <= sub_wire82(30);
	sub_wire2(175, 31)    <= sub_wire82(31);
	sub_wire2(175, 32)    <= sub_wire82(32);
	sub_wire2(175, 33)    <= sub_wire82(33);
	sub_wire2(175, 34)    <= sub_wire82(34);
	sub_wire2(175, 35)    <= sub_wire82(35);
	sub_wire2(175, 36)    <= sub_wire82(36);
	sub_wire2(175, 37)    <= sub_wire82(37);
	sub_wire2(175, 38)    <= sub_wire82(38);
	sub_wire2(175, 39)    <= sub_wire82(39);
	sub_wire2(174, 0)    <= sub_wire83(0);
	sub_wire2(174, 1)    <= sub_wire83(1);
	sub_wire2(174, 2)    <= sub_wire83(2);
	sub_wire2(174, 3)    <= sub_wire83(3);
	sub_wire2(174, 4)    <= sub_wire83(4);
	sub_wire2(174, 5)    <= sub_wire83(5);
	sub_wire2(174, 6)    <= sub_wire83(6);
	sub_wire2(174, 7)    <= sub_wire83(7);
	sub_wire2(174, 8)    <= sub_wire83(8);
	sub_wire2(174, 9)    <= sub_wire83(9);
	sub_wire2(174, 10)    <= sub_wire83(10);
	sub_wire2(174, 11)    <= sub_wire83(11);
	sub_wire2(174, 12)    <= sub_wire83(12);
	sub_wire2(174, 13)    <= sub_wire83(13);
	sub_wire2(174, 14)    <= sub_wire83(14);
	sub_wire2(174, 15)    <= sub_wire83(15);
	sub_wire2(174, 16)    <= sub_wire83(16);
	sub_wire2(174, 17)    <= sub_wire83(17);
	sub_wire2(174, 18)    <= sub_wire83(18);
	sub_wire2(174, 19)    <= sub_wire83(19);
	sub_wire2(174, 20)    <= sub_wire83(20);
	sub_wire2(174, 21)    <= sub_wire83(21);
	sub_wire2(174, 22)    <= sub_wire83(22);
	sub_wire2(174, 23)    <= sub_wire83(23);
	sub_wire2(174, 24)    <= sub_wire83(24);
	sub_wire2(174, 25)    <= sub_wire83(25);
	sub_wire2(174, 26)    <= sub_wire83(26);
	sub_wire2(174, 27)    <= sub_wire83(27);
	sub_wire2(174, 28)    <= sub_wire83(28);
	sub_wire2(174, 29)    <= sub_wire83(29);
	sub_wire2(174, 30)    <= sub_wire83(30);
	sub_wire2(174, 31)    <= sub_wire83(31);
	sub_wire2(174, 32)    <= sub_wire83(32);
	sub_wire2(174, 33)    <= sub_wire83(33);
	sub_wire2(174, 34)    <= sub_wire83(34);
	sub_wire2(174, 35)    <= sub_wire83(35);
	sub_wire2(174, 36)    <= sub_wire83(36);
	sub_wire2(174, 37)    <= sub_wire83(37);
	sub_wire2(174, 38)    <= sub_wire83(38);
	sub_wire2(174, 39)    <= sub_wire83(39);
	sub_wire2(173, 0)    <= sub_wire84(0);
	sub_wire2(173, 1)    <= sub_wire84(1);
	sub_wire2(173, 2)    <= sub_wire84(2);
	sub_wire2(173, 3)    <= sub_wire84(3);
	sub_wire2(173, 4)    <= sub_wire84(4);
	sub_wire2(173, 5)    <= sub_wire84(5);
	sub_wire2(173, 6)    <= sub_wire84(6);
	sub_wire2(173, 7)    <= sub_wire84(7);
	sub_wire2(173, 8)    <= sub_wire84(8);
	sub_wire2(173, 9)    <= sub_wire84(9);
	sub_wire2(173, 10)    <= sub_wire84(10);
	sub_wire2(173, 11)    <= sub_wire84(11);
	sub_wire2(173, 12)    <= sub_wire84(12);
	sub_wire2(173, 13)    <= sub_wire84(13);
	sub_wire2(173, 14)    <= sub_wire84(14);
	sub_wire2(173, 15)    <= sub_wire84(15);
	sub_wire2(173, 16)    <= sub_wire84(16);
	sub_wire2(173, 17)    <= sub_wire84(17);
	sub_wire2(173, 18)    <= sub_wire84(18);
	sub_wire2(173, 19)    <= sub_wire84(19);
	sub_wire2(173, 20)    <= sub_wire84(20);
	sub_wire2(173, 21)    <= sub_wire84(21);
	sub_wire2(173, 22)    <= sub_wire84(22);
	sub_wire2(173, 23)    <= sub_wire84(23);
	sub_wire2(173, 24)    <= sub_wire84(24);
	sub_wire2(173, 25)    <= sub_wire84(25);
	sub_wire2(173, 26)    <= sub_wire84(26);
	sub_wire2(173, 27)    <= sub_wire84(27);
	sub_wire2(173, 28)    <= sub_wire84(28);
	sub_wire2(173, 29)    <= sub_wire84(29);
	sub_wire2(173, 30)    <= sub_wire84(30);
	sub_wire2(173, 31)    <= sub_wire84(31);
	sub_wire2(173, 32)    <= sub_wire84(32);
	sub_wire2(173, 33)    <= sub_wire84(33);
	sub_wire2(173, 34)    <= sub_wire84(34);
	sub_wire2(173, 35)    <= sub_wire84(35);
	sub_wire2(173, 36)    <= sub_wire84(36);
	sub_wire2(173, 37)    <= sub_wire84(37);
	sub_wire2(173, 38)    <= sub_wire84(38);
	sub_wire2(173, 39)    <= sub_wire84(39);
	sub_wire2(172, 0)    <= sub_wire85(0);
	sub_wire2(172, 1)    <= sub_wire85(1);
	sub_wire2(172, 2)    <= sub_wire85(2);
	sub_wire2(172, 3)    <= sub_wire85(3);
	sub_wire2(172, 4)    <= sub_wire85(4);
	sub_wire2(172, 5)    <= sub_wire85(5);
	sub_wire2(172, 6)    <= sub_wire85(6);
	sub_wire2(172, 7)    <= sub_wire85(7);
	sub_wire2(172, 8)    <= sub_wire85(8);
	sub_wire2(172, 9)    <= sub_wire85(9);
	sub_wire2(172, 10)    <= sub_wire85(10);
	sub_wire2(172, 11)    <= sub_wire85(11);
	sub_wire2(172, 12)    <= sub_wire85(12);
	sub_wire2(172, 13)    <= sub_wire85(13);
	sub_wire2(172, 14)    <= sub_wire85(14);
	sub_wire2(172, 15)    <= sub_wire85(15);
	sub_wire2(172, 16)    <= sub_wire85(16);
	sub_wire2(172, 17)    <= sub_wire85(17);
	sub_wire2(172, 18)    <= sub_wire85(18);
	sub_wire2(172, 19)    <= sub_wire85(19);
	sub_wire2(172, 20)    <= sub_wire85(20);
	sub_wire2(172, 21)    <= sub_wire85(21);
	sub_wire2(172, 22)    <= sub_wire85(22);
	sub_wire2(172, 23)    <= sub_wire85(23);
	sub_wire2(172, 24)    <= sub_wire85(24);
	sub_wire2(172, 25)    <= sub_wire85(25);
	sub_wire2(172, 26)    <= sub_wire85(26);
	sub_wire2(172, 27)    <= sub_wire85(27);
	sub_wire2(172, 28)    <= sub_wire85(28);
	sub_wire2(172, 29)    <= sub_wire85(29);
	sub_wire2(172, 30)    <= sub_wire85(30);
	sub_wire2(172, 31)    <= sub_wire85(31);
	sub_wire2(172, 32)    <= sub_wire85(32);
	sub_wire2(172, 33)    <= sub_wire85(33);
	sub_wire2(172, 34)    <= sub_wire85(34);
	sub_wire2(172, 35)    <= sub_wire85(35);
	sub_wire2(172, 36)    <= sub_wire85(36);
	sub_wire2(172, 37)    <= sub_wire85(37);
	sub_wire2(172, 38)    <= sub_wire85(38);
	sub_wire2(172, 39)    <= sub_wire85(39);
	sub_wire2(171, 0)    <= sub_wire86(0);
	sub_wire2(171, 1)    <= sub_wire86(1);
	sub_wire2(171, 2)    <= sub_wire86(2);
	sub_wire2(171, 3)    <= sub_wire86(3);
	sub_wire2(171, 4)    <= sub_wire86(4);
	sub_wire2(171, 5)    <= sub_wire86(5);
	sub_wire2(171, 6)    <= sub_wire86(6);
	sub_wire2(171, 7)    <= sub_wire86(7);
	sub_wire2(171, 8)    <= sub_wire86(8);
	sub_wire2(171, 9)    <= sub_wire86(9);
	sub_wire2(171, 10)    <= sub_wire86(10);
	sub_wire2(171, 11)    <= sub_wire86(11);
	sub_wire2(171, 12)    <= sub_wire86(12);
	sub_wire2(171, 13)    <= sub_wire86(13);
	sub_wire2(171, 14)    <= sub_wire86(14);
	sub_wire2(171, 15)    <= sub_wire86(15);
	sub_wire2(171, 16)    <= sub_wire86(16);
	sub_wire2(171, 17)    <= sub_wire86(17);
	sub_wire2(171, 18)    <= sub_wire86(18);
	sub_wire2(171, 19)    <= sub_wire86(19);
	sub_wire2(171, 20)    <= sub_wire86(20);
	sub_wire2(171, 21)    <= sub_wire86(21);
	sub_wire2(171, 22)    <= sub_wire86(22);
	sub_wire2(171, 23)    <= sub_wire86(23);
	sub_wire2(171, 24)    <= sub_wire86(24);
	sub_wire2(171, 25)    <= sub_wire86(25);
	sub_wire2(171, 26)    <= sub_wire86(26);
	sub_wire2(171, 27)    <= sub_wire86(27);
	sub_wire2(171, 28)    <= sub_wire86(28);
	sub_wire2(171, 29)    <= sub_wire86(29);
	sub_wire2(171, 30)    <= sub_wire86(30);
	sub_wire2(171, 31)    <= sub_wire86(31);
	sub_wire2(171, 32)    <= sub_wire86(32);
	sub_wire2(171, 33)    <= sub_wire86(33);
	sub_wire2(171, 34)    <= sub_wire86(34);
	sub_wire2(171, 35)    <= sub_wire86(35);
	sub_wire2(171, 36)    <= sub_wire86(36);
	sub_wire2(171, 37)    <= sub_wire86(37);
	sub_wire2(171, 38)    <= sub_wire86(38);
	sub_wire2(171, 39)    <= sub_wire86(39);
	sub_wire2(170, 0)    <= sub_wire87(0);
	sub_wire2(170, 1)    <= sub_wire87(1);
	sub_wire2(170, 2)    <= sub_wire87(2);
	sub_wire2(170, 3)    <= sub_wire87(3);
	sub_wire2(170, 4)    <= sub_wire87(4);
	sub_wire2(170, 5)    <= sub_wire87(5);
	sub_wire2(170, 6)    <= sub_wire87(6);
	sub_wire2(170, 7)    <= sub_wire87(7);
	sub_wire2(170, 8)    <= sub_wire87(8);
	sub_wire2(170, 9)    <= sub_wire87(9);
	sub_wire2(170, 10)    <= sub_wire87(10);
	sub_wire2(170, 11)    <= sub_wire87(11);
	sub_wire2(170, 12)    <= sub_wire87(12);
	sub_wire2(170, 13)    <= sub_wire87(13);
	sub_wire2(170, 14)    <= sub_wire87(14);
	sub_wire2(170, 15)    <= sub_wire87(15);
	sub_wire2(170, 16)    <= sub_wire87(16);
	sub_wire2(170, 17)    <= sub_wire87(17);
	sub_wire2(170, 18)    <= sub_wire87(18);
	sub_wire2(170, 19)    <= sub_wire87(19);
	sub_wire2(170, 20)    <= sub_wire87(20);
	sub_wire2(170, 21)    <= sub_wire87(21);
	sub_wire2(170, 22)    <= sub_wire87(22);
	sub_wire2(170, 23)    <= sub_wire87(23);
	sub_wire2(170, 24)    <= sub_wire87(24);
	sub_wire2(170, 25)    <= sub_wire87(25);
	sub_wire2(170, 26)    <= sub_wire87(26);
	sub_wire2(170, 27)    <= sub_wire87(27);
	sub_wire2(170, 28)    <= sub_wire87(28);
	sub_wire2(170, 29)    <= sub_wire87(29);
	sub_wire2(170, 30)    <= sub_wire87(30);
	sub_wire2(170, 31)    <= sub_wire87(31);
	sub_wire2(170, 32)    <= sub_wire87(32);
	sub_wire2(170, 33)    <= sub_wire87(33);
	sub_wire2(170, 34)    <= sub_wire87(34);
	sub_wire2(170, 35)    <= sub_wire87(35);
	sub_wire2(170, 36)    <= sub_wire87(36);
	sub_wire2(170, 37)    <= sub_wire87(37);
	sub_wire2(170, 38)    <= sub_wire87(38);
	sub_wire2(170, 39)    <= sub_wire87(39);
	sub_wire2(169, 0)    <= sub_wire88(0);
	sub_wire2(169, 1)    <= sub_wire88(1);
	sub_wire2(169, 2)    <= sub_wire88(2);
	sub_wire2(169, 3)    <= sub_wire88(3);
	sub_wire2(169, 4)    <= sub_wire88(4);
	sub_wire2(169, 5)    <= sub_wire88(5);
	sub_wire2(169, 6)    <= sub_wire88(6);
	sub_wire2(169, 7)    <= sub_wire88(7);
	sub_wire2(169, 8)    <= sub_wire88(8);
	sub_wire2(169, 9)    <= sub_wire88(9);
	sub_wire2(169, 10)    <= sub_wire88(10);
	sub_wire2(169, 11)    <= sub_wire88(11);
	sub_wire2(169, 12)    <= sub_wire88(12);
	sub_wire2(169, 13)    <= sub_wire88(13);
	sub_wire2(169, 14)    <= sub_wire88(14);
	sub_wire2(169, 15)    <= sub_wire88(15);
	sub_wire2(169, 16)    <= sub_wire88(16);
	sub_wire2(169, 17)    <= sub_wire88(17);
	sub_wire2(169, 18)    <= sub_wire88(18);
	sub_wire2(169, 19)    <= sub_wire88(19);
	sub_wire2(169, 20)    <= sub_wire88(20);
	sub_wire2(169, 21)    <= sub_wire88(21);
	sub_wire2(169, 22)    <= sub_wire88(22);
	sub_wire2(169, 23)    <= sub_wire88(23);
	sub_wire2(169, 24)    <= sub_wire88(24);
	sub_wire2(169, 25)    <= sub_wire88(25);
	sub_wire2(169, 26)    <= sub_wire88(26);
	sub_wire2(169, 27)    <= sub_wire88(27);
	sub_wire2(169, 28)    <= sub_wire88(28);
	sub_wire2(169, 29)    <= sub_wire88(29);
	sub_wire2(169, 30)    <= sub_wire88(30);
	sub_wire2(169, 31)    <= sub_wire88(31);
	sub_wire2(169, 32)    <= sub_wire88(32);
	sub_wire2(169, 33)    <= sub_wire88(33);
	sub_wire2(169, 34)    <= sub_wire88(34);
	sub_wire2(169, 35)    <= sub_wire88(35);
	sub_wire2(169, 36)    <= sub_wire88(36);
	sub_wire2(169, 37)    <= sub_wire88(37);
	sub_wire2(169, 38)    <= sub_wire88(38);
	sub_wire2(169, 39)    <= sub_wire88(39);
	sub_wire2(168, 0)    <= sub_wire89(0);
	sub_wire2(168, 1)    <= sub_wire89(1);
	sub_wire2(168, 2)    <= sub_wire89(2);
	sub_wire2(168, 3)    <= sub_wire89(3);
	sub_wire2(168, 4)    <= sub_wire89(4);
	sub_wire2(168, 5)    <= sub_wire89(5);
	sub_wire2(168, 6)    <= sub_wire89(6);
	sub_wire2(168, 7)    <= sub_wire89(7);
	sub_wire2(168, 8)    <= sub_wire89(8);
	sub_wire2(168, 9)    <= sub_wire89(9);
	sub_wire2(168, 10)    <= sub_wire89(10);
	sub_wire2(168, 11)    <= sub_wire89(11);
	sub_wire2(168, 12)    <= sub_wire89(12);
	sub_wire2(168, 13)    <= sub_wire89(13);
	sub_wire2(168, 14)    <= sub_wire89(14);
	sub_wire2(168, 15)    <= sub_wire89(15);
	sub_wire2(168, 16)    <= sub_wire89(16);
	sub_wire2(168, 17)    <= sub_wire89(17);
	sub_wire2(168, 18)    <= sub_wire89(18);
	sub_wire2(168, 19)    <= sub_wire89(19);
	sub_wire2(168, 20)    <= sub_wire89(20);
	sub_wire2(168, 21)    <= sub_wire89(21);
	sub_wire2(168, 22)    <= sub_wire89(22);
	sub_wire2(168, 23)    <= sub_wire89(23);
	sub_wire2(168, 24)    <= sub_wire89(24);
	sub_wire2(168, 25)    <= sub_wire89(25);
	sub_wire2(168, 26)    <= sub_wire89(26);
	sub_wire2(168, 27)    <= sub_wire89(27);
	sub_wire2(168, 28)    <= sub_wire89(28);
	sub_wire2(168, 29)    <= sub_wire89(29);
	sub_wire2(168, 30)    <= sub_wire89(30);
	sub_wire2(168, 31)    <= sub_wire89(31);
	sub_wire2(168, 32)    <= sub_wire89(32);
	sub_wire2(168, 33)    <= sub_wire89(33);
	sub_wire2(168, 34)    <= sub_wire89(34);
	sub_wire2(168, 35)    <= sub_wire89(35);
	sub_wire2(168, 36)    <= sub_wire89(36);
	sub_wire2(168, 37)    <= sub_wire89(37);
	sub_wire2(168, 38)    <= sub_wire89(38);
	sub_wire2(168, 39)    <= sub_wire89(39);
	sub_wire2(167, 0)    <= sub_wire90(0);
	sub_wire2(167, 1)    <= sub_wire90(1);
	sub_wire2(167, 2)    <= sub_wire90(2);
	sub_wire2(167, 3)    <= sub_wire90(3);
	sub_wire2(167, 4)    <= sub_wire90(4);
	sub_wire2(167, 5)    <= sub_wire90(5);
	sub_wire2(167, 6)    <= sub_wire90(6);
	sub_wire2(167, 7)    <= sub_wire90(7);
	sub_wire2(167, 8)    <= sub_wire90(8);
	sub_wire2(167, 9)    <= sub_wire90(9);
	sub_wire2(167, 10)    <= sub_wire90(10);
	sub_wire2(167, 11)    <= sub_wire90(11);
	sub_wire2(167, 12)    <= sub_wire90(12);
	sub_wire2(167, 13)    <= sub_wire90(13);
	sub_wire2(167, 14)    <= sub_wire90(14);
	sub_wire2(167, 15)    <= sub_wire90(15);
	sub_wire2(167, 16)    <= sub_wire90(16);
	sub_wire2(167, 17)    <= sub_wire90(17);
	sub_wire2(167, 18)    <= sub_wire90(18);
	sub_wire2(167, 19)    <= sub_wire90(19);
	sub_wire2(167, 20)    <= sub_wire90(20);
	sub_wire2(167, 21)    <= sub_wire90(21);
	sub_wire2(167, 22)    <= sub_wire90(22);
	sub_wire2(167, 23)    <= sub_wire90(23);
	sub_wire2(167, 24)    <= sub_wire90(24);
	sub_wire2(167, 25)    <= sub_wire90(25);
	sub_wire2(167, 26)    <= sub_wire90(26);
	sub_wire2(167, 27)    <= sub_wire90(27);
	sub_wire2(167, 28)    <= sub_wire90(28);
	sub_wire2(167, 29)    <= sub_wire90(29);
	sub_wire2(167, 30)    <= sub_wire90(30);
	sub_wire2(167, 31)    <= sub_wire90(31);
	sub_wire2(167, 32)    <= sub_wire90(32);
	sub_wire2(167, 33)    <= sub_wire90(33);
	sub_wire2(167, 34)    <= sub_wire90(34);
	sub_wire2(167, 35)    <= sub_wire90(35);
	sub_wire2(167, 36)    <= sub_wire90(36);
	sub_wire2(167, 37)    <= sub_wire90(37);
	sub_wire2(167, 38)    <= sub_wire90(38);
	sub_wire2(167, 39)    <= sub_wire90(39);
	sub_wire2(166, 0)    <= sub_wire91(0);
	sub_wire2(166, 1)    <= sub_wire91(1);
	sub_wire2(166, 2)    <= sub_wire91(2);
	sub_wire2(166, 3)    <= sub_wire91(3);
	sub_wire2(166, 4)    <= sub_wire91(4);
	sub_wire2(166, 5)    <= sub_wire91(5);
	sub_wire2(166, 6)    <= sub_wire91(6);
	sub_wire2(166, 7)    <= sub_wire91(7);
	sub_wire2(166, 8)    <= sub_wire91(8);
	sub_wire2(166, 9)    <= sub_wire91(9);
	sub_wire2(166, 10)    <= sub_wire91(10);
	sub_wire2(166, 11)    <= sub_wire91(11);
	sub_wire2(166, 12)    <= sub_wire91(12);
	sub_wire2(166, 13)    <= sub_wire91(13);
	sub_wire2(166, 14)    <= sub_wire91(14);
	sub_wire2(166, 15)    <= sub_wire91(15);
	sub_wire2(166, 16)    <= sub_wire91(16);
	sub_wire2(166, 17)    <= sub_wire91(17);
	sub_wire2(166, 18)    <= sub_wire91(18);
	sub_wire2(166, 19)    <= sub_wire91(19);
	sub_wire2(166, 20)    <= sub_wire91(20);
	sub_wire2(166, 21)    <= sub_wire91(21);
	sub_wire2(166, 22)    <= sub_wire91(22);
	sub_wire2(166, 23)    <= sub_wire91(23);
	sub_wire2(166, 24)    <= sub_wire91(24);
	sub_wire2(166, 25)    <= sub_wire91(25);
	sub_wire2(166, 26)    <= sub_wire91(26);
	sub_wire2(166, 27)    <= sub_wire91(27);
	sub_wire2(166, 28)    <= sub_wire91(28);
	sub_wire2(166, 29)    <= sub_wire91(29);
	sub_wire2(166, 30)    <= sub_wire91(30);
	sub_wire2(166, 31)    <= sub_wire91(31);
	sub_wire2(166, 32)    <= sub_wire91(32);
	sub_wire2(166, 33)    <= sub_wire91(33);
	sub_wire2(166, 34)    <= sub_wire91(34);
	sub_wire2(166, 35)    <= sub_wire91(35);
	sub_wire2(166, 36)    <= sub_wire91(36);
	sub_wire2(166, 37)    <= sub_wire91(37);
	sub_wire2(166, 38)    <= sub_wire91(38);
	sub_wire2(166, 39)    <= sub_wire91(39);
	sub_wire2(165, 0)    <= sub_wire92(0);
	sub_wire2(165, 1)    <= sub_wire92(1);
	sub_wire2(165, 2)    <= sub_wire92(2);
	sub_wire2(165, 3)    <= sub_wire92(3);
	sub_wire2(165, 4)    <= sub_wire92(4);
	sub_wire2(165, 5)    <= sub_wire92(5);
	sub_wire2(165, 6)    <= sub_wire92(6);
	sub_wire2(165, 7)    <= sub_wire92(7);
	sub_wire2(165, 8)    <= sub_wire92(8);
	sub_wire2(165, 9)    <= sub_wire92(9);
	sub_wire2(165, 10)    <= sub_wire92(10);
	sub_wire2(165, 11)    <= sub_wire92(11);
	sub_wire2(165, 12)    <= sub_wire92(12);
	sub_wire2(165, 13)    <= sub_wire92(13);
	sub_wire2(165, 14)    <= sub_wire92(14);
	sub_wire2(165, 15)    <= sub_wire92(15);
	sub_wire2(165, 16)    <= sub_wire92(16);
	sub_wire2(165, 17)    <= sub_wire92(17);
	sub_wire2(165, 18)    <= sub_wire92(18);
	sub_wire2(165, 19)    <= sub_wire92(19);
	sub_wire2(165, 20)    <= sub_wire92(20);
	sub_wire2(165, 21)    <= sub_wire92(21);
	sub_wire2(165, 22)    <= sub_wire92(22);
	sub_wire2(165, 23)    <= sub_wire92(23);
	sub_wire2(165, 24)    <= sub_wire92(24);
	sub_wire2(165, 25)    <= sub_wire92(25);
	sub_wire2(165, 26)    <= sub_wire92(26);
	sub_wire2(165, 27)    <= sub_wire92(27);
	sub_wire2(165, 28)    <= sub_wire92(28);
	sub_wire2(165, 29)    <= sub_wire92(29);
	sub_wire2(165, 30)    <= sub_wire92(30);
	sub_wire2(165, 31)    <= sub_wire92(31);
	sub_wire2(165, 32)    <= sub_wire92(32);
	sub_wire2(165, 33)    <= sub_wire92(33);
	sub_wire2(165, 34)    <= sub_wire92(34);
	sub_wire2(165, 35)    <= sub_wire92(35);
	sub_wire2(165, 36)    <= sub_wire92(36);
	sub_wire2(165, 37)    <= sub_wire92(37);
	sub_wire2(165, 38)    <= sub_wire92(38);
	sub_wire2(165, 39)    <= sub_wire92(39);
	sub_wire2(164, 0)    <= sub_wire93(0);
	sub_wire2(164, 1)    <= sub_wire93(1);
	sub_wire2(164, 2)    <= sub_wire93(2);
	sub_wire2(164, 3)    <= sub_wire93(3);
	sub_wire2(164, 4)    <= sub_wire93(4);
	sub_wire2(164, 5)    <= sub_wire93(5);
	sub_wire2(164, 6)    <= sub_wire93(6);
	sub_wire2(164, 7)    <= sub_wire93(7);
	sub_wire2(164, 8)    <= sub_wire93(8);
	sub_wire2(164, 9)    <= sub_wire93(9);
	sub_wire2(164, 10)    <= sub_wire93(10);
	sub_wire2(164, 11)    <= sub_wire93(11);
	sub_wire2(164, 12)    <= sub_wire93(12);
	sub_wire2(164, 13)    <= sub_wire93(13);
	sub_wire2(164, 14)    <= sub_wire93(14);
	sub_wire2(164, 15)    <= sub_wire93(15);
	sub_wire2(164, 16)    <= sub_wire93(16);
	sub_wire2(164, 17)    <= sub_wire93(17);
	sub_wire2(164, 18)    <= sub_wire93(18);
	sub_wire2(164, 19)    <= sub_wire93(19);
	sub_wire2(164, 20)    <= sub_wire93(20);
	sub_wire2(164, 21)    <= sub_wire93(21);
	sub_wire2(164, 22)    <= sub_wire93(22);
	sub_wire2(164, 23)    <= sub_wire93(23);
	sub_wire2(164, 24)    <= sub_wire93(24);
	sub_wire2(164, 25)    <= sub_wire93(25);
	sub_wire2(164, 26)    <= sub_wire93(26);
	sub_wire2(164, 27)    <= sub_wire93(27);
	sub_wire2(164, 28)    <= sub_wire93(28);
	sub_wire2(164, 29)    <= sub_wire93(29);
	sub_wire2(164, 30)    <= sub_wire93(30);
	sub_wire2(164, 31)    <= sub_wire93(31);
	sub_wire2(164, 32)    <= sub_wire93(32);
	sub_wire2(164, 33)    <= sub_wire93(33);
	sub_wire2(164, 34)    <= sub_wire93(34);
	sub_wire2(164, 35)    <= sub_wire93(35);
	sub_wire2(164, 36)    <= sub_wire93(36);
	sub_wire2(164, 37)    <= sub_wire93(37);
	sub_wire2(164, 38)    <= sub_wire93(38);
	sub_wire2(164, 39)    <= sub_wire93(39);
	sub_wire2(163, 0)    <= sub_wire94(0);
	sub_wire2(163, 1)    <= sub_wire94(1);
	sub_wire2(163, 2)    <= sub_wire94(2);
	sub_wire2(163, 3)    <= sub_wire94(3);
	sub_wire2(163, 4)    <= sub_wire94(4);
	sub_wire2(163, 5)    <= sub_wire94(5);
	sub_wire2(163, 6)    <= sub_wire94(6);
	sub_wire2(163, 7)    <= sub_wire94(7);
	sub_wire2(163, 8)    <= sub_wire94(8);
	sub_wire2(163, 9)    <= sub_wire94(9);
	sub_wire2(163, 10)    <= sub_wire94(10);
	sub_wire2(163, 11)    <= sub_wire94(11);
	sub_wire2(163, 12)    <= sub_wire94(12);
	sub_wire2(163, 13)    <= sub_wire94(13);
	sub_wire2(163, 14)    <= sub_wire94(14);
	sub_wire2(163, 15)    <= sub_wire94(15);
	sub_wire2(163, 16)    <= sub_wire94(16);
	sub_wire2(163, 17)    <= sub_wire94(17);
	sub_wire2(163, 18)    <= sub_wire94(18);
	sub_wire2(163, 19)    <= sub_wire94(19);
	sub_wire2(163, 20)    <= sub_wire94(20);
	sub_wire2(163, 21)    <= sub_wire94(21);
	sub_wire2(163, 22)    <= sub_wire94(22);
	sub_wire2(163, 23)    <= sub_wire94(23);
	sub_wire2(163, 24)    <= sub_wire94(24);
	sub_wire2(163, 25)    <= sub_wire94(25);
	sub_wire2(163, 26)    <= sub_wire94(26);
	sub_wire2(163, 27)    <= sub_wire94(27);
	sub_wire2(163, 28)    <= sub_wire94(28);
	sub_wire2(163, 29)    <= sub_wire94(29);
	sub_wire2(163, 30)    <= sub_wire94(30);
	sub_wire2(163, 31)    <= sub_wire94(31);
	sub_wire2(163, 32)    <= sub_wire94(32);
	sub_wire2(163, 33)    <= sub_wire94(33);
	sub_wire2(163, 34)    <= sub_wire94(34);
	sub_wire2(163, 35)    <= sub_wire94(35);
	sub_wire2(163, 36)    <= sub_wire94(36);
	sub_wire2(163, 37)    <= sub_wire94(37);
	sub_wire2(163, 38)    <= sub_wire94(38);
	sub_wire2(163, 39)    <= sub_wire94(39);
	sub_wire2(162, 0)    <= sub_wire95(0);
	sub_wire2(162, 1)    <= sub_wire95(1);
	sub_wire2(162, 2)    <= sub_wire95(2);
	sub_wire2(162, 3)    <= sub_wire95(3);
	sub_wire2(162, 4)    <= sub_wire95(4);
	sub_wire2(162, 5)    <= sub_wire95(5);
	sub_wire2(162, 6)    <= sub_wire95(6);
	sub_wire2(162, 7)    <= sub_wire95(7);
	sub_wire2(162, 8)    <= sub_wire95(8);
	sub_wire2(162, 9)    <= sub_wire95(9);
	sub_wire2(162, 10)    <= sub_wire95(10);
	sub_wire2(162, 11)    <= sub_wire95(11);
	sub_wire2(162, 12)    <= sub_wire95(12);
	sub_wire2(162, 13)    <= sub_wire95(13);
	sub_wire2(162, 14)    <= sub_wire95(14);
	sub_wire2(162, 15)    <= sub_wire95(15);
	sub_wire2(162, 16)    <= sub_wire95(16);
	sub_wire2(162, 17)    <= sub_wire95(17);
	sub_wire2(162, 18)    <= sub_wire95(18);
	sub_wire2(162, 19)    <= sub_wire95(19);
	sub_wire2(162, 20)    <= sub_wire95(20);
	sub_wire2(162, 21)    <= sub_wire95(21);
	sub_wire2(162, 22)    <= sub_wire95(22);
	sub_wire2(162, 23)    <= sub_wire95(23);
	sub_wire2(162, 24)    <= sub_wire95(24);
	sub_wire2(162, 25)    <= sub_wire95(25);
	sub_wire2(162, 26)    <= sub_wire95(26);
	sub_wire2(162, 27)    <= sub_wire95(27);
	sub_wire2(162, 28)    <= sub_wire95(28);
	sub_wire2(162, 29)    <= sub_wire95(29);
	sub_wire2(162, 30)    <= sub_wire95(30);
	sub_wire2(162, 31)    <= sub_wire95(31);
	sub_wire2(162, 32)    <= sub_wire95(32);
	sub_wire2(162, 33)    <= sub_wire95(33);
	sub_wire2(162, 34)    <= sub_wire95(34);
	sub_wire2(162, 35)    <= sub_wire95(35);
	sub_wire2(162, 36)    <= sub_wire95(36);
	sub_wire2(162, 37)    <= sub_wire95(37);
	sub_wire2(162, 38)    <= sub_wire95(38);
	sub_wire2(162, 39)    <= sub_wire95(39);
	sub_wire2(161, 0)    <= sub_wire96(0);
	sub_wire2(161, 1)    <= sub_wire96(1);
	sub_wire2(161, 2)    <= sub_wire96(2);
	sub_wire2(161, 3)    <= sub_wire96(3);
	sub_wire2(161, 4)    <= sub_wire96(4);
	sub_wire2(161, 5)    <= sub_wire96(5);
	sub_wire2(161, 6)    <= sub_wire96(6);
	sub_wire2(161, 7)    <= sub_wire96(7);
	sub_wire2(161, 8)    <= sub_wire96(8);
	sub_wire2(161, 9)    <= sub_wire96(9);
	sub_wire2(161, 10)    <= sub_wire96(10);
	sub_wire2(161, 11)    <= sub_wire96(11);
	sub_wire2(161, 12)    <= sub_wire96(12);
	sub_wire2(161, 13)    <= sub_wire96(13);
	sub_wire2(161, 14)    <= sub_wire96(14);
	sub_wire2(161, 15)    <= sub_wire96(15);
	sub_wire2(161, 16)    <= sub_wire96(16);
	sub_wire2(161, 17)    <= sub_wire96(17);
	sub_wire2(161, 18)    <= sub_wire96(18);
	sub_wire2(161, 19)    <= sub_wire96(19);
	sub_wire2(161, 20)    <= sub_wire96(20);
	sub_wire2(161, 21)    <= sub_wire96(21);
	sub_wire2(161, 22)    <= sub_wire96(22);
	sub_wire2(161, 23)    <= sub_wire96(23);
	sub_wire2(161, 24)    <= sub_wire96(24);
	sub_wire2(161, 25)    <= sub_wire96(25);
	sub_wire2(161, 26)    <= sub_wire96(26);
	sub_wire2(161, 27)    <= sub_wire96(27);
	sub_wire2(161, 28)    <= sub_wire96(28);
	sub_wire2(161, 29)    <= sub_wire96(29);
	sub_wire2(161, 30)    <= sub_wire96(30);
	sub_wire2(161, 31)    <= sub_wire96(31);
	sub_wire2(161, 32)    <= sub_wire96(32);
	sub_wire2(161, 33)    <= sub_wire96(33);
	sub_wire2(161, 34)    <= sub_wire96(34);
	sub_wire2(161, 35)    <= sub_wire96(35);
	sub_wire2(161, 36)    <= sub_wire96(36);
	sub_wire2(161, 37)    <= sub_wire96(37);
	sub_wire2(161, 38)    <= sub_wire96(38);
	sub_wire2(161, 39)    <= sub_wire96(39);
	sub_wire2(160, 0)    <= sub_wire97(0);
	sub_wire2(160, 1)    <= sub_wire97(1);
	sub_wire2(160, 2)    <= sub_wire97(2);
	sub_wire2(160, 3)    <= sub_wire97(3);
	sub_wire2(160, 4)    <= sub_wire97(4);
	sub_wire2(160, 5)    <= sub_wire97(5);
	sub_wire2(160, 6)    <= sub_wire97(6);
	sub_wire2(160, 7)    <= sub_wire97(7);
	sub_wire2(160, 8)    <= sub_wire97(8);
	sub_wire2(160, 9)    <= sub_wire97(9);
	sub_wire2(160, 10)    <= sub_wire97(10);
	sub_wire2(160, 11)    <= sub_wire97(11);
	sub_wire2(160, 12)    <= sub_wire97(12);
	sub_wire2(160, 13)    <= sub_wire97(13);
	sub_wire2(160, 14)    <= sub_wire97(14);
	sub_wire2(160, 15)    <= sub_wire97(15);
	sub_wire2(160, 16)    <= sub_wire97(16);
	sub_wire2(160, 17)    <= sub_wire97(17);
	sub_wire2(160, 18)    <= sub_wire97(18);
	sub_wire2(160, 19)    <= sub_wire97(19);
	sub_wire2(160, 20)    <= sub_wire97(20);
	sub_wire2(160, 21)    <= sub_wire97(21);
	sub_wire2(160, 22)    <= sub_wire97(22);
	sub_wire2(160, 23)    <= sub_wire97(23);
	sub_wire2(160, 24)    <= sub_wire97(24);
	sub_wire2(160, 25)    <= sub_wire97(25);
	sub_wire2(160, 26)    <= sub_wire97(26);
	sub_wire2(160, 27)    <= sub_wire97(27);
	sub_wire2(160, 28)    <= sub_wire97(28);
	sub_wire2(160, 29)    <= sub_wire97(29);
	sub_wire2(160, 30)    <= sub_wire97(30);
	sub_wire2(160, 31)    <= sub_wire97(31);
	sub_wire2(160, 32)    <= sub_wire97(32);
	sub_wire2(160, 33)    <= sub_wire97(33);
	sub_wire2(160, 34)    <= sub_wire97(34);
	sub_wire2(160, 35)    <= sub_wire97(35);
	sub_wire2(160, 36)    <= sub_wire97(36);
	sub_wire2(160, 37)    <= sub_wire97(37);
	sub_wire2(160, 38)    <= sub_wire97(38);
	sub_wire2(160, 39)    <= sub_wire97(39);
	sub_wire2(159, 0)    <= sub_wire98(0);
	sub_wire2(159, 1)    <= sub_wire98(1);
	sub_wire2(159, 2)    <= sub_wire98(2);
	sub_wire2(159, 3)    <= sub_wire98(3);
	sub_wire2(159, 4)    <= sub_wire98(4);
	sub_wire2(159, 5)    <= sub_wire98(5);
	sub_wire2(159, 6)    <= sub_wire98(6);
	sub_wire2(159, 7)    <= sub_wire98(7);
	sub_wire2(159, 8)    <= sub_wire98(8);
	sub_wire2(159, 9)    <= sub_wire98(9);
	sub_wire2(159, 10)    <= sub_wire98(10);
	sub_wire2(159, 11)    <= sub_wire98(11);
	sub_wire2(159, 12)    <= sub_wire98(12);
	sub_wire2(159, 13)    <= sub_wire98(13);
	sub_wire2(159, 14)    <= sub_wire98(14);
	sub_wire2(159, 15)    <= sub_wire98(15);
	sub_wire2(159, 16)    <= sub_wire98(16);
	sub_wire2(159, 17)    <= sub_wire98(17);
	sub_wire2(159, 18)    <= sub_wire98(18);
	sub_wire2(159, 19)    <= sub_wire98(19);
	sub_wire2(159, 20)    <= sub_wire98(20);
	sub_wire2(159, 21)    <= sub_wire98(21);
	sub_wire2(159, 22)    <= sub_wire98(22);
	sub_wire2(159, 23)    <= sub_wire98(23);
	sub_wire2(159, 24)    <= sub_wire98(24);
	sub_wire2(159, 25)    <= sub_wire98(25);
	sub_wire2(159, 26)    <= sub_wire98(26);
	sub_wire2(159, 27)    <= sub_wire98(27);
	sub_wire2(159, 28)    <= sub_wire98(28);
	sub_wire2(159, 29)    <= sub_wire98(29);
	sub_wire2(159, 30)    <= sub_wire98(30);
	sub_wire2(159, 31)    <= sub_wire98(31);
	sub_wire2(159, 32)    <= sub_wire98(32);
	sub_wire2(159, 33)    <= sub_wire98(33);
	sub_wire2(159, 34)    <= sub_wire98(34);
	sub_wire2(159, 35)    <= sub_wire98(35);
	sub_wire2(159, 36)    <= sub_wire98(36);
	sub_wire2(159, 37)    <= sub_wire98(37);
	sub_wire2(159, 38)    <= sub_wire98(38);
	sub_wire2(159, 39)    <= sub_wire98(39);
	sub_wire2(158, 0)    <= sub_wire99(0);
	sub_wire2(158, 1)    <= sub_wire99(1);
	sub_wire2(158, 2)    <= sub_wire99(2);
	sub_wire2(158, 3)    <= sub_wire99(3);
	sub_wire2(158, 4)    <= sub_wire99(4);
	sub_wire2(158, 5)    <= sub_wire99(5);
	sub_wire2(158, 6)    <= sub_wire99(6);
	sub_wire2(158, 7)    <= sub_wire99(7);
	sub_wire2(158, 8)    <= sub_wire99(8);
	sub_wire2(158, 9)    <= sub_wire99(9);
	sub_wire2(158, 10)    <= sub_wire99(10);
	sub_wire2(158, 11)    <= sub_wire99(11);
	sub_wire2(158, 12)    <= sub_wire99(12);
	sub_wire2(158, 13)    <= sub_wire99(13);
	sub_wire2(158, 14)    <= sub_wire99(14);
	sub_wire2(158, 15)    <= sub_wire99(15);
	sub_wire2(158, 16)    <= sub_wire99(16);
	sub_wire2(158, 17)    <= sub_wire99(17);
	sub_wire2(158, 18)    <= sub_wire99(18);
	sub_wire2(158, 19)    <= sub_wire99(19);
	sub_wire2(158, 20)    <= sub_wire99(20);
	sub_wire2(158, 21)    <= sub_wire99(21);
	sub_wire2(158, 22)    <= sub_wire99(22);
	sub_wire2(158, 23)    <= sub_wire99(23);
	sub_wire2(158, 24)    <= sub_wire99(24);
	sub_wire2(158, 25)    <= sub_wire99(25);
	sub_wire2(158, 26)    <= sub_wire99(26);
	sub_wire2(158, 27)    <= sub_wire99(27);
	sub_wire2(158, 28)    <= sub_wire99(28);
	sub_wire2(158, 29)    <= sub_wire99(29);
	sub_wire2(158, 30)    <= sub_wire99(30);
	sub_wire2(158, 31)    <= sub_wire99(31);
	sub_wire2(158, 32)    <= sub_wire99(32);
	sub_wire2(158, 33)    <= sub_wire99(33);
	sub_wire2(158, 34)    <= sub_wire99(34);
	sub_wire2(158, 35)    <= sub_wire99(35);
	sub_wire2(158, 36)    <= sub_wire99(36);
	sub_wire2(158, 37)    <= sub_wire99(37);
	sub_wire2(158, 38)    <= sub_wire99(38);
	sub_wire2(158, 39)    <= sub_wire99(39);
	sub_wire2(157, 0)    <= sub_wire100(0);
	sub_wire2(157, 1)    <= sub_wire100(1);
	sub_wire2(157, 2)    <= sub_wire100(2);
	sub_wire2(157, 3)    <= sub_wire100(3);
	sub_wire2(157, 4)    <= sub_wire100(4);
	sub_wire2(157, 5)    <= sub_wire100(5);
	sub_wire2(157, 6)    <= sub_wire100(6);
	sub_wire2(157, 7)    <= sub_wire100(7);
	sub_wire2(157, 8)    <= sub_wire100(8);
	sub_wire2(157, 9)    <= sub_wire100(9);
	sub_wire2(157, 10)    <= sub_wire100(10);
	sub_wire2(157, 11)    <= sub_wire100(11);
	sub_wire2(157, 12)    <= sub_wire100(12);
	sub_wire2(157, 13)    <= sub_wire100(13);
	sub_wire2(157, 14)    <= sub_wire100(14);
	sub_wire2(157, 15)    <= sub_wire100(15);
	sub_wire2(157, 16)    <= sub_wire100(16);
	sub_wire2(157, 17)    <= sub_wire100(17);
	sub_wire2(157, 18)    <= sub_wire100(18);
	sub_wire2(157, 19)    <= sub_wire100(19);
	sub_wire2(157, 20)    <= sub_wire100(20);
	sub_wire2(157, 21)    <= sub_wire100(21);
	sub_wire2(157, 22)    <= sub_wire100(22);
	sub_wire2(157, 23)    <= sub_wire100(23);
	sub_wire2(157, 24)    <= sub_wire100(24);
	sub_wire2(157, 25)    <= sub_wire100(25);
	sub_wire2(157, 26)    <= sub_wire100(26);
	sub_wire2(157, 27)    <= sub_wire100(27);
	sub_wire2(157, 28)    <= sub_wire100(28);
	sub_wire2(157, 29)    <= sub_wire100(29);
	sub_wire2(157, 30)    <= sub_wire100(30);
	sub_wire2(157, 31)    <= sub_wire100(31);
	sub_wire2(157, 32)    <= sub_wire100(32);
	sub_wire2(157, 33)    <= sub_wire100(33);
	sub_wire2(157, 34)    <= sub_wire100(34);
	sub_wire2(157, 35)    <= sub_wire100(35);
	sub_wire2(157, 36)    <= sub_wire100(36);
	sub_wire2(157, 37)    <= sub_wire100(37);
	sub_wire2(157, 38)    <= sub_wire100(38);
	sub_wire2(157, 39)    <= sub_wire100(39);
	sub_wire2(156, 0)    <= sub_wire101(0);
	sub_wire2(156, 1)    <= sub_wire101(1);
	sub_wire2(156, 2)    <= sub_wire101(2);
	sub_wire2(156, 3)    <= sub_wire101(3);
	sub_wire2(156, 4)    <= sub_wire101(4);
	sub_wire2(156, 5)    <= sub_wire101(5);
	sub_wire2(156, 6)    <= sub_wire101(6);
	sub_wire2(156, 7)    <= sub_wire101(7);
	sub_wire2(156, 8)    <= sub_wire101(8);
	sub_wire2(156, 9)    <= sub_wire101(9);
	sub_wire2(156, 10)    <= sub_wire101(10);
	sub_wire2(156, 11)    <= sub_wire101(11);
	sub_wire2(156, 12)    <= sub_wire101(12);
	sub_wire2(156, 13)    <= sub_wire101(13);
	sub_wire2(156, 14)    <= sub_wire101(14);
	sub_wire2(156, 15)    <= sub_wire101(15);
	sub_wire2(156, 16)    <= sub_wire101(16);
	sub_wire2(156, 17)    <= sub_wire101(17);
	sub_wire2(156, 18)    <= sub_wire101(18);
	sub_wire2(156, 19)    <= sub_wire101(19);
	sub_wire2(156, 20)    <= sub_wire101(20);
	sub_wire2(156, 21)    <= sub_wire101(21);
	sub_wire2(156, 22)    <= sub_wire101(22);
	sub_wire2(156, 23)    <= sub_wire101(23);
	sub_wire2(156, 24)    <= sub_wire101(24);
	sub_wire2(156, 25)    <= sub_wire101(25);
	sub_wire2(156, 26)    <= sub_wire101(26);
	sub_wire2(156, 27)    <= sub_wire101(27);
	sub_wire2(156, 28)    <= sub_wire101(28);
	sub_wire2(156, 29)    <= sub_wire101(29);
	sub_wire2(156, 30)    <= sub_wire101(30);
	sub_wire2(156, 31)    <= sub_wire101(31);
	sub_wire2(156, 32)    <= sub_wire101(32);
	sub_wire2(156, 33)    <= sub_wire101(33);
	sub_wire2(156, 34)    <= sub_wire101(34);
	sub_wire2(156, 35)    <= sub_wire101(35);
	sub_wire2(156, 36)    <= sub_wire101(36);
	sub_wire2(156, 37)    <= sub_wire101(37);
	sub_wire2(156, 38)    <= sub_wire101(38);
	sub_wire2(156, 39)    <= sub_wire101(39);
	sub_wire2(155, 0)    <= sub_wire102(0);
	sub_wire2(155, 1)    <= sub_wire102(1);
	sub_wire2(155, 2)    <= sub_wire102(2);
	sub_wire2(155, 3)    <= sub_wire102(3);
	sub_wire2(155, 4)    <= sub_wire102(4);
	sub_wire2(155, 5)    <= sub_wire102(5);
	sub_wire2(155, 6)    <= sub_wire102(6);
	sub_wire2(155, 7)    <= sub_wire102(7);
	sub_wire2(155, 8)    <= sub_wire102(8);
	sub_wire2(155, 9)    <= sub_wire102(9);
	sub_wire2(155, 10)    <= sub_wire102(10);
	sub_wire2(155, 11)    <= sub_wire102(11);
	sub_wire2(155, 12)    <= sub_wire102(12);
	sub_wire2(155, 13)    <= sub_wire102(13);
	sub_wire2(155, 14)    <= sub_wire102(14);
	sub_wire2(155, 15)    <= sub_wire102(15);
	sub_wire2(155, 16)    <= sub_wire102(16);
	sub_wire2(155, 17)    <= sub_wire102(17);
	sub_wire2(155, 18)    <= sub_wire102(18);
	sub_wire2(155, 19)    <= sub_wire102(19);
	sub_wire2(155, 20)    <= sub_wire102(20);
	sub_wire2(155, 21)    <= sub_wire102(21);
	sub_wire2(155, 22)    <= sub_wire102(22);
	sub_wire2(155, 23)    <= sub_wire102(23);
	sub_wire2(155, 24)    <= sub_wire102(24);
	sub_wire2(155, 25)    <= sub_wire102(25);
	sub_wire2(155, 26)    <= sub_wire102(26);
	sub_wire2(155, 27)    <= sub_wire102(27);
	sub_wire2(155, 28)    <= sub_wire102(28);
	sub_wire2(155, 29)    <= sub_wire102(29);
	sub_wire2(155, 30)    <= sub_wire102(30);
	sub_wire2(155, 31)    <= sub_wire102(31);
	sub_wire2(155, 32)    <= sub_wire102(32);
	sub_wire2(155, 33)    <= sub_wire102(33);
	sub_wire2(155, 34)    <= sub_wire102(34);
	sub_wire2(155, 35)    <= sub_wire102(35);
	sub_wire2(155, 36)    <= sub_wire102(36);
	sub_wire2(155, 37)    <= sub_wire102(37);
	sub_wire2(155, 38)    <= sub_wire102(38);
	sub_wire2(155, 39)    <= sub_wire102(39);
	sub_wire2(154, 0)    <= sub_wire103(0);
	sub_wire2(154, 1)    <= sub_wire103(1);
	sub_wire2(154, 2)    <= sub_wire103(2);
	sub_wire2(154, 3)    <= sub_wire103(3);
	sub_wire2(154, 4)    <= sub_wire103(4);
	sub_wire2(154, 5)    <= sub_wire103(5);
	sub_wire2(154, 6)    <= sub_wire103(6);
	sub_wire2(154, 7)    <= sub_wire103(7);
	sub_wire2(154, 8)    <= sub_wire103(8);
	sub_wire2(154, 9)    <= sub_wire103(9);
	sub_wire2(154, 10)    <= sub_wire103(10);
	sub_wire2(154, 11)    <= sub_wire103(11);
	sub_wire2(154, 12)    <= sub_wire103(12);
	sub_wire2(154, 13)    <= sub_wire103(13);
	sub_wire2(154, 14)    <= sub_wire103(14);
	sub_wire2(154, 15)    <= sub_wire103(15);
	sub_wire2(154, 16)    <= sub_wire103(16);
	sub_wire2(154, 17)    <= sub_wire103(17);
	sub_wire2(154, 18)    <= sub_wire103(18);
	sub_wire2(154, 19)    <= sub_wire103(19);
	sub_wire2(154, 20)    <= sub_wire103(20);
	sub_wire2(154, 21)    <= sub_wire103(21);
	sub_wire2(154, 22)    <= sub_wire103(22);
	sub_wire2(154, 23)    <= sub_wire103(23);
	sub_wire2(154, 24)    <= sub_wire103(24);
	sub_wire2(154, 25)    <= sub_wire103(25);
	sub_wire2(154, 26)    <= sub_wire103(26);
	sub_wire2(154, 27)    <= sub_wire103(27);
	sub_wire2(154, 28)    <= sub_wire103(28);
	sub_wire2(154, 29)    <= sub_wire103(29);
	sub_wire2(154, 30)    <= sub_wire103(30);
	sub_wire2(154, 31)    <= sub_wire103(31);
	sub_wire2(154, 32)    <= sub_wire103(32);
	sub_wire2(154, 33)    <= sub_wire103(33);
	sub_wire2(154, 34)    <= sub_wire103(34);
	sub_wire2(154, 35)    <= sub_wire103(35);
	sub_wire2(154, 36)    <= sub_wire103(36);
	sub_wire2(154, 37)    <= sub_wire103(37);
	sub_wire2(154, 38)    <= sub_wire103(38);
	sub_wire2(154, 39)    <= sub_wire103(39);
	sub_wire2(153, 0)    <= sub_wire104(0);
	sub_wire2(153, 1)    <= sub_wire104(1);
	sub_wire2(153, 2)    <= sub_wire104(2);
	sub_wire2(153, 3)    <= sub_wire104(3);
	sub_wire2(153, 4)    <= sub_wire104(4);
	sub_wire2(153, 5)    <= sub_wire104(5);
	sub_wire2(153, 6)    <= sub_wire104(6);
	sub_wire2(153, 7)    <= sub_wire104(7);
	sub_wire2(153, 8)    <= sub_wire104(8);
	sub_wire2(153, 9)    <= sub_wire104(9);
	sub_wire2(153, 10)    <= sub_wire104(10);
	sub_wire2(153, 11)    <= sub_wire104(11);
	sub_wire2(153, 12)    <= sub_wire104(12);
	sub_wire2(153, 13)    <= sub_wire104(13);
	sub_wire2(153, 14)    <= sub_wire104(14);
	sub_wire2(153, 15)    <= sub_wire104(15);
	sub_wire2(153, 16)    <= sub_wire104(16);
	sub_wire2(153, 17)    <= sub_wire104(17);
	sub_wire2(153, 18)    <= sub_wire104(18);
	sub_wire2(153, 19)    <= sub_wire104(19);
	sub_wire2(153, 20)    <= sub_wire104(20);
	sub_wire2(153, 21)    <= sub_wire104(21);
	sub_wire2(153, 22)    <= sub_wire104(22);
	sub_wire2(153, 23)    <= sub_wire104(23);
	sub_wire2(153, 24)    <= sub_wire104(24);
	sub_wire2(153, 25)    <= sub_wire104(25);
	sub_wire2(153, 26)    <= sub_wire104(26);
	sub_wire2(153, 27)    <= sub_wire104(27);
	sub_wire2(153, 28)    <= sub_wire104(28);
	sub_wire2(153, 29)    <= sub_wire104(29);
	sub_wire2(153, 30)    <= sub_wire104(30);
	sub_wire2(153, 31)    <= sub_wire104(31);
	sub_wire2(153, 32)    <= sub_wire104(32);
	sub_wire2(153, 33)    <= sub_wire104(33);
	sub_wire2(153, 34)    <= sub_wire104(34);
	sub_wire2(153, 35)    <= sub_wire104(35);
	sub_wire2(153, 36)    <= sub_wire104(36);
	sub_wire2(153, 37)    <= sub_wire104(37);
	sub_wire2(153, 38)    <= sub_wire104(38);
	sub_wire2(153, 39)    <= sub_wire104(39);
	sub_wire2(152, 0)    <= sub_wire105(0);
	sub_wire2(152, 1)    <= sub_wire105(1);
	sub_wire2(152, 2)    <= sub_wire105(2);
	sub_wire2(152, 3)    <= sub_wire105(3);
	sub_wire2(152, 4)    <= sub_wire105(4);
	sub_wire2(152, 5)    <= sub_wire105(5);
	sub_wire2(152, 6)    <= sub_wire105(6);
	sub_wire2(152, 7)    <= sub_wire105(7);
	sub_wire2(152, 8)    <= sub_wire105(8);
	sub_wire2(152, 9)    <= sub_wire105(9);
	sub_wire2(152, 10)    <= sub_wire105(10);
	sub_wire2(152, 11)    <= sub_wire105(11);
	sub_wire2(152, 12)    <= sub_wire105(12);
	sub_wire2(152, 13)    <= sub_wire105(13);
	sub_wire2(152, 14)    <= sub_wire105(14);
	sub_wire2(152, 15)    <= sub_wire105(15);
	sub_wire2(152, 16)    <= sub_wire105(16);
	sub_wire2(152, 17)    <= sub_wire105(17);
	sub_wire2(152, 18)    <= sub_wire105(18);
	sub_wire2(152, 19)    <= sub_wire105(19);
	sub_wire2(152, 20)    <= sub_wire105(20);
	sub_wire2(152, 21)    <= sub_wire105(21);
	sub_wire2(152, 22)    <= sub_wire105(22);
	sub_wire2(152, 23)    <= sub_wire105(23);
	sub_wire2(152, 24)    <= sub_wire105(24);
	sub_wire2(152, 25)    <= sub_wire105(25);
	sub_wire2(152, 26)    <= sub_wire105(26);
	sub_wire2(152, 27)    <= sub_wire105(27);
	sub_wire2(152, 28)    <= sub_wire105(28);
	sub_wire2(152, 29)    <= sub_wire105(29);
	sub_wire2(152, 30)    <= sub_wire105(30);
	sub_wire2(152, 31)    <= sub_wire105(31);
	sub_wire2(152, 32)    <= sub_wire105(32);
	sub_wire2(152, 33)    <= sub_wire105(33);
	sub_wire2(152, 34)    <= sub_wire105(34);
	sub_wire2(152, 35)    <= sub_wire105(35);
	sub_wire2(152, 36)    <= sub_wire105(36);
	sub_wire2(152, 37)    <= sub_wire105(37);
	sub_wire2(152, 38)    <= sub_wire105(38);
	sub_wire2(152, 39)    <= sub_wire105(39);
	sub_wire2(151, 0)    <= sub_wire106(0);
	sub_wire2(151, 1)    <= sub_wire106(1);
	sub_wire2(151, 2)    <= sub_wire106(2);
	sub_wire2(151, 3)    <= sub_wire106(3);
	sub_wire2(151, 4)    <= sub_wire106(4);
	sub_wire2(151, 5)    <= sub_wire106(5);
	sub_wire2(151, 6)    <= sub_wire106(6);
	sub_wire2(151, 7)    <= sub_wire106(7);
	sub_wire2(151, 8)    <= sub_wire106(8);
	sub_wire2(151, 9)    <= sub_wire106(9);
	sub_wire2(151, 10)    <= sub_wire106(10);
	sub_wire2(151, 11)    <= sub_wire106(11);
	sub_wire2(151, 12)    <= sub_wire106(12);
	sub_wire2(151, 13)    <= sub_wire106(13);
	sub_wire2(151, 14)    <= sub_wire106(14);
	sub_wire2(151, 15)    <= sub_wire106(15);
	sub_wire2(151, 16)    <= sub_wire106(16);
	sub_wire2(151, 17)    <= sub_wire106(17);
	sub_wire2(151, 18)    <= sub_wire106(18);
	sub_wire2(151, 19)    <= sub_wire106(19);
	sub_wire2(151, 20)    <= sub_wire106(20);
	sub_wire2(151, 21)    <= sub_wire106(21);
	sub_wire2(151, 22)    <= sub_wire106(22);
	sub_wire2(151, 23)    <= sub_wire106(23);
	sub_wire2(151, 24)    <= sub_wire106(24);
	sub_wire2(151, 25)    <= sub_wire106(25);
	sub_wire2(151, 26)    <= sub_wire106(26);
	sub_wire2(151, 27)    <= sub_wire106(27);
	sub_wire2(151, 28)    <= sub_wire106(28);
	sub_wire2(151, 29)    <= sub_wire106(29);
	sub_wire2(151, 30)    <= sub_wire106(30);
	sub_wire2(151, 31)    <= sub_wire106(31);
	sub_wire2(151, 32)    <= sub_wire106(32);
	sub_wire2(151, 33)    <= sub_wire106(33);
	sub_wire2(151, 34)    <= sub_wire106(34);
	sub_wire2(151, 35)    <= sub_wire106(35);
	sub_wire2(151, 36)    <= sub_wire106(36);
	sub_wire2(151, 37)    <= sub_wire106(37);
	sub_wire2(151, 38)    <= sub_wire106(38);
	sub_wire2(151, 39)    <= sub_wire106(39);
	sub_wire2(150, 0)    <= sub_wire107(0);
	sub_wire2(150, 1)    <= sub_wire107(1);
	sub_wire2(150, 2)    <= sub_wire107(2);
	sub_wire2(150, 3)    <= sub_wire107(3);
	sub_wire2(150, 4)    <= sub_wire107(4);
	sub_wire2(150, 5)    <= sub_wire107(5);
	sub_wire2(150, 6)    <= sub_wire107(6);
	sub_wire2(150, 7)    <= sub_wire107(7);
	sub_wire2(150, 8)    <= sub_wire107(8);
	sub_wire2(150, 9)    <= sub_wire107(9);
	sub_wire2(150, 10)    <= sub_wire107(10);
	sub_wire2(150, 11)    <= sub_wire107(11);
	sub_wire2(150, 12)    <= sub_wire107(12);
	sub_wire2(150, 13)    <= sub_wire107(13);
	sub_wire2(150, 14)    <= sub_wire107(14);
	sub_wire2(150, 15)    <= sub_wire107(15);
	sub_wire2(150, 16)    <= sub_wire107(16);
	sub_wire2(150, 17)    <= sub_wire107(17);
	sub_wire2(150, 18)    <= sub_wire107(18);
	sub_wire2(150, 19)    <= sub_wire107(19);
	sub_wire2(150, 20)    <= sub_wire107(20);
	sub_wire2(150, 21)    <= sub_wire107(21);
	sub_wire2(150, 22)    <= sub_wire107(22);
	sub_wire2(150, 23)    <= sub_wire107(23);
	sub_wire2(150, 24)    <= sub_wire107(24);
	sub_wire2(150, 25)    <= sub_wire107(25);
	sub_wire2(150, 26)    <= sub_wire107(26);
	sub_wire2(150, 27)    <= sub_wire107(27);
	sub_wire2(150, 28)    <= sub_wire107(28);
	sub_wire2(150, 29)    <= sub_wire107(29);
	sub_wire2(150, 30)    <= sub_wire107(30);
	sub_wire2(150, 31)    <= sub_wire107(31);
	sub_wire2(150, 32)    <= sub_wire107(32);
	sub_wire2(150, 33)    <= sub_wire107(33);
	sub_wire2(150, 34)    <= sub_wire107(34);
	sub_wire2(150, 35)    <= sub_wire107(35);
	sub_wire2(150, 36)    <= sub_wire107(36);
	sub_wire2(150, 37)    <= sub_wire107(37);
	sub_wire2(150, 38)    <= sub_wire107(38);
	sub_wire2(150, 39)    <= sub_wire107(39);
	sub_wire2(149, 0)    <= sub_wire108(0);
	sub_wire2(149, 1)    <= sub_wire108(1);
	sub_wire2(149, 2)    <= sub_wire108(2);
	sub_wire2(149, 3)    <= sub_wire108(3);
	sub_wire2(149, 4)    <= sub_wire108(4);
	sub_wire2(149, 5)    <= sub_wire108(5);
	sub_wire2(149, 6)    <= sub_wire108(6);
	sub_wire2(149, 7)    <= sub_wire108(7);
	sub_wire2(149, 8)    <= sub_wire108(8);
	sub_wire2(149, 9)    <= sub_wire108(9);
	sub_wire2(149, 10)    <= sub_wire108(10);
	sub_wire2(149, 11)    <= sub_wire108(11);
	sub_wire2(149, 12)    <= sub_wire108(12);
	sub_wire2(149, 13)    <= sub_wire108(13);
	sub_wire2(149, 14)    <= sub_wire108(14);
	sub_wire2(149, 15)    <= sub_wire108(15);
	sub_wire2(149, 16)    <= sub_wire108(16);
	sub_wire2(149, 17)    <= sub_wire108(17);
	sub_wire2(149, 18)    <= sub_wire108(18);
	sub_wire2(149, 19)    <= sub_wire108(19);
	sub_wire2(149, 20)    <= sub_wire108(20);
	sub_wire2(149, 21)    <= sub_wire108(21);
	sub_wire2(149, 22)    <= sub_wire108(22);
	sub_wire2(149, 23)    <= sub_wire108(23);
	sub_wire2(149, 24)    <= sub_wire108(24);
	sub_wire2(149, 25)    <= sub_wire108(25);
	sub_wire2(149, 26)    <= sub_wire108(26);
	sub_wire2(149, 27)    <= sub_wire108(27);
	sub_wire2(149, 28)    <= sub_wire108(28);
	sub_wire2(149, 29)    <= sub_wire108(29);
	sub_wire2(149, 30)    <= sub_wire108(30);
	sub_wire2(149, 31)    <= sub_wire108(31);
	sub_wire2(149, 32)    <= sub_wire108(32);
	sub_wire2(149, 33)    <= sub_wire108(33);
	sub_wire2(149, 34)    <= sub_wire108(34);
	sub_wire2(149, 35)    <= sub_wire108(35);
	sub_wire2(149, 36)    <= sub_wire108(36);
	sub_wire2(149, 37)    <= sub_wire108(37);
	sub_wire2(149, 38)    <= sub_wire108(38);
	sub_wire2(149, 39)    <= sub_wire108(39);
	sub_wire2(148, 0)    <= sub_wire109(0);
	sub_wire2(148, 1)    <= sub_wire109(1);
	sub_wire2(148, 2)    <= sub_wire109(2);
	sub_wire2(148, 3)    <= sub_wire109(3);
	sub_wire2(148, 4)    <= sub_wire109(4);
	sub_wire2(148, 5)    <= sub_wire109(5);
	sub_wire2(148, 6)    <= sub_wire109(6);
	sub_wire2(148, 7)    <= sub_wire109(7);
	sub_wire2(148, 8)    <= sub_wire109(8);
	sub_wire2(148, 9)    <= sub_wire109(9);
	sub_wire2(148, 10)    <= sub_wire109(10);
	sub_wire2(148, 11)    <= sub_wire109(11);
	sub_wire2(148, 12)    <= sub_wire109(12);
	sub_wire2(148, 13)    <= sub_wire109(13);
	sub_wire2(148, 14)    <= sub_wire109(14);
	sub_wire2(148, 15)    <= sub_wire109(15);
	sub_wire2(148, 16)    <= sub_wire109(16);
	sub_wire2(148, 17)    <= sub_wire109(17);
	sub_wire2(148, 18)    <= sub_wire109(18);
	sub_wire2(148, 19)    <= sub_wire109(19);
	sub_wire2(148, 20)    <= sub_wire109(20);
	sub_wire2(148, 21)    <= sub_wire109(21);
	sub_wire2(148, 22)    <= sub_wire109(22);
	sub_wire2(148, 23)    <= sub_wire109(23);
	sub_wire2(148, 24)    <= sub_wire109(24);
	sub_wire2(148, 25)    <= sub_wire109(25);
	sub_wire2(148, 26)    <= sub_wire109(26);
	sub_wire2(148, 27)    <= sub_wire109(27);
	sub_wire2(148, 28)    <= sub_wire109(28);
	sub_wire2(148, 29)    <= sub_wire109(29);
	sub_wire2(148, 30)    <= sub_wire109(30);
	sub_wire2(148, 31)    <= sub_wire109(31);
	sub_wire2(148, 32)    <= sub_wire109(32);
	sub_wire2(148, 33)    <= sub_wire109(33);
	sub_wire2(148, 34)    <= sub_wire109(34);
	sub_wire2(148, 35)    <= sub_wire109(35);
	sub_wire2(148, 36)    <= sub_wire109(36);
	sub_wire2(148, 37)    <= sub_wire109(37);
	sub_wire2(148, 38)    <= sub_wire109(38);
	sub_wire2(148, 39)    <= sub_wire109(39);
	sub_wire2(147, 0)    <= sub_wire110(0);
	sub_wire2(147, 1)    <= sub_wire110(1);
	sub_wire2(147, 2)    <= sub_wire110(2);
	sub_wire2(147, 3)    <= sub_wire110(3);
	sub_wire2(147, 4)    <= sub_wire110(4);
	sub_wire2(147, 5)    <= sub_wire110(5);
	sub_wire2(147, 6)    <= sub_wire110(6);
	sub_wire2(147, 7)    <= sub_wire110(7);
	sub_wire2(147, 8)    <= sub_wire110(8);
	sub_wire2(147, 9)    <= sub_wire110(9);
	sub_wire2(147, 10)    <= sub_wire110(10);
	sub_wire2(147, 11)    <= sub_wire110(11);
	sub_wire2(147, 12)    <= sub_wire110(12);
	sub_wire2(147, 13)    <= sub_wire110(13);
	sub_wire2(147, 14)    <= sub_wire110(14);
	sub_wire2(147, 15)    <= sub_wire110(15);
	sub_wire2(147, 16)    <= sub_wire110(16);
	sub_wire2(147, 17)    <= sub_wire110(17);
	sub_wire2(147, 18)    <= sub_wire110(18);
	sub_wire2(147, 19)    <= sub_wire110(19);
	sub_wire2(147, 20)    <= sub_wire110(20);
	sub_wire2(147, 21)    <= sub_wire110(21);
	sub_wire2(147, 22)    <= sub_wire110(22);
	sub_wire2(147, 23)    <= sub_wire110(23);
	sub_wire2(147, 24)    <= sub_wire110(24);
	sub_wire2(147, 25)    <= sub_wire110(25);
	sub_wire2(147, 26)    <= sub_wire110(26);
	sub_wire2(147, 27)    <= sub_wire110(27);
	sub_wire2(147, 28)    <= sub_wire110(28);
	sub_wire2(147, 29)    <= sub_wire110(29);
	sub_wire2(147, 30)    <= sub_wire110(30);
	sub_wire2(147, 31)    <= sub_wire110(31);
	sub_wire2(147, 32)    <= sub_wire110(32);
	sub_wire2(147, 33)    <= sub_wire110(33);
	sub_wire2(147, 34)    <= sub_wire110(34);
	sub_wire2(147, 35)    <= sub_wire110(35);
	sub_wire2(147, 36)    <= sub_wire110(36);
	sub_wire2(147, 37)    <= sub_wire110(37);
	sub_wire2(147, 38)    <= sub_wire110(38);
	sub_wire2(147, 39)    <= sub_wire110(39);
	sub_wire2(146, 0)    <= sub_wire111(0);
	sub_wire2(146, 1)    <= sub_wire111(1);
	sub_wire2(146, 2)    <= sub_wire111(2);
	sub_wire2(146, 3)    <= sub_wire111(3);
	sub_wire2(146, 4)    <= sub_wire111(4);
	sub_wire2(146, 5)    <= sub_wire111(5);
	sub_wire2(146, 6)    <= sub_wire111(6);
	sub_wire2(146, 7)    <= sub_wire111(7);
	sub_wire2(146, 8)    <= sub_wire111(8);
	sub_wire2(146, 9)    <= sub_wire111(9);
	sub_wire2(146, 10)    <= sub_wire111(10);
	sub_wire2(146, 11)    <= sub_wire111(11);
	sub_wire2(146, 12)    <= sub_wire111(12);
	sub_wire2(146, 13)    <= sub_wire111(13);
	sub_wire2(146, 14)    <= sub_wire111(14);
	sub_wire2(146, 15)    <= sub_wire111(15);
	sub_wire2(146, 16)    <= sub_wire111(16);
	sub_wire2(146, 17)    <= sub_wire111(17);
	sub_wire2(146, 18)    <= sub_wire111(18);
	sub_wire2(146, 19)    <= sub_wire111(19);
	sub_wire2(146, 20)    <= sub_wire111(20);
	sub_wire2(146, 21)    <= sub_wire111(21);
	sub_wire2(146, 22)    <= sub_wire111(22);
	sub_wire2(146, 23)    <= sub_wire111(23);
	sub_wire2(146, 24)    <= sub_wire111(24);
	sub_wire2(146, 25)    <= sub_wire111(25);
	sub_wire2(146, 26)    <= sub_wire111(26);
	sub_wire2(146, 27)    <= sub_wire111(27);
	sub_wire2(146, 28)    <= sub_wire111(28);
	sub_wire2(146, 29)    <= sub_wire111(29);
	sub_wire2(146, 30)    <= sub_wire111(30);
	sub_wire2(146, 31)    <= sub_wire111(31);
	sub_wire2(146, 32)    <= sub_wire111(32);
	sub_wire2(146, 33)    <= sub_wire111(33);
	sub_wire2(146, 34)    <= sub_wire111(34);
	sub_wire2(146, 35)    <= sub_wire111(35);
	sub_wire2(146, 36)    <= sub_wire111(36);
	sub_wire2(146, 37)    <= sub_wire111(37);
	sub_wire2(146, 38)    <= sub_wire111(38);
	sub_wire2(146, 39)    <= sub_wire111(39);
	sub_wire2(145, 0)    <= sub_wire112(0);
	sub_wire2(145, 1)    <= sub_wire112(1);
	sub_wire2(145, 2)    <= sub_wire112(2);
	sub_wire2(145, 3)    <= sub_wire112(3);
	sub_wire2(145, 4)    <= sub_wire112(4);
	sub_wire2(145, 5)    <= sub_wire112(5);
	sub_wire2(145, 6)    <= sub_wire112(6);
	sub_wire2(145, 7)    <= sub_wire112(7);
	sub_wire2(145, 8)    <= sub_wire112(8);
	sub_wire2(145, 9)    <= sub_wire112(9);
	sub_wire2(145, 10)    <= sub_wire112(10);
	sub_wire2(145, 11)    <= sub_wire112(11);
	sub_wire2(145, 12)    <= sub_wire112(12);
	sub_wire2(145, 13)    <= sub_wire112(13);
	sub_wire2(145, 14)    <= sub_wire112(14);
	sub_wire2(145, 15)    <= sub_wire112(15);
	sub_wire2(145, 16)    <= sub_wire112(16);
	sub_wire2(145, 17)    <= sub_wire112(17);
	sub_wire2(145, 18)    <= sub_wire112(18);
	sub_wire2(145, 19)    <= sub_wire112(19);
	sub_wire2(145, 20)    <= sub_wire112(20);
	sub_wire2(145, 21)    <= sub_wire112(21);
	sub_wire2(145, 22)    <= sub_wire112(22);
	sub_wire2(145, 23)    <= sub_wire112(23);
	sub_wire2(145, 24)    <= sub_wire112(24);
	sub_wire2(145, 25)    <= sub_wire112(25);
	sub_wire2(145, 26)    <= sub_wire112(26);
	sub_wire2(145, 27)    <= sub_wire112(27);
	sub_wire2(145, 28)    <= sub_wire112(28);
	sub_wire2(145, 29)    <= sub_wire112(29);
	sub_wire2(145, 30)    <= sub_wire112(30);
	sub_wire2(145, 31)    <= sub_wire112(31);
	sub_wire2(145, 32)    <= sub_wire112(32);
	sub_wire2(145, 33)    <= sub_wire112(33);
	sub_wire2(145, 34)    <= sub_wire112(34);
	sub_wire2(145, 35)    <= sub_wire112(35);
	sub_wire2(145, 36)    <= sub_wire112(36);
	sub_wire2(145, 37)    <= sub_wire112(37);
	sub_wire2(145, 38)    <= sub_wire112(38);
	sub_wire2(145, 39)    <= sub_wire112(39);
	sub_wire2(144, 0)    <= sub_wire113(0);
	sub_wire2(144, 1)    <= sub_wire113(1);
	sub_wire2(144, 2)    <= sub_wire113(2);
	sub_wire2(144, 3)    <= sub_wire113(3);
	sub_wire2(144, 4)    <= sub_wire113(4);
	sub_wire2(144, 5)    <= sub_wire113(5);
	sub_wire2(144, 6)    <= sub_wire113(6);
	sub_wire2(144, 7)    <= sub_wire113(7);
	sub_wire2(144, 8)    <= sub_wire113(8);
	sub_wire2(144, 9)    <= sub_wire113(9);
	sub_wire2(144, 10)    <= sub_wire113(10);
	sub_wire2(144, 11)    <= sub_wire113(11);
	sub_wire2(144, 12)    <= sub_wire113(12);
	sub_wire2(144, 13)    <= sub_wire113(13);
	sub_wire2(144, 14)    <= sub_wire113(14);
	sub_wire2(144, 15)    <= sub_wire113(15);
	sub_wire2(144, 16)    <= sub_wire113(16);
	sub_wire2(144, 17)    <= sub_wire113(17);
	sub_wire2(144, 18)    <= sub_wire113(18);
	sub_wire2(144, 19)    <= sub_wire113(19);
	sub_wire2(144, 20)    <= sub_wire113(20);
	sub_wire2(144, 21)    <= sub_wire113(21);
	sub_wire2(144, 22)    <= sub_wire113(22);
	sub_wire2(144, 23)    <= sub_wire113(23);
	sub_wire2(144, 24)    <= sub_wire113(24);
	sub_wire2(144, 25)    <= sub_wire113(25);
	sub_wire2(144, 26)    <= sub_wire113(26);
	sub_wire2(144, 27)    <= sub_wire113(27);
	sub_wire2(144, 28)    <= sub_wire113(28);
	sub_wire2(144, 29)    <= sub_wire113(29);
	sub_wire2(144, 30)    <= sub_wire113(30);
	sub_wire2(144, 31)    <= sub_wire113(31);
	sub_wire2(144, 32)    <= sub_wire113(32);
	sub_wire2(144, 33)    <= sub_wire113(33);
	sub_wire2(144, 34)    <= sub_wire113(34);
	sub_wire2(144, 35)    <= sub_wire113(35);
	sub_wire2(144, 36)    <= sub_wire113(36);
	sub_wire2(144, 37)    <= sub_wire113(37);
	sub_wire2(144, 38)    <= sub_wire113(38);
	sub_wire2(144, 39)    <= sub_wire113(39);
	sub_wire2(143, 0)    <= sub_wire114(0);
	sub_wire2(143, 1)    <= sub_wire114(1);
	sub_wire2(143, 2)    <= sub_wire114(2);
	sub_wire2(143, 3)    <= sub_wire114(3);
	sub_wire2(143, 4)    <= sub_wire114(4);
	sub_wire2(143, 5)    <= sub_wire114(5);
	sub_wire2(143, 6)    <= sub_wire114(6);
	sub_wire2(143, 7)    <= sub_wire114(7);
	sub_wire2(143, 8)    <= sub_wire114(8);
	sub_wire2(143, 9)    <= sub_wire114(9);
	sub_wire2(143, 10)    <= sub_wire114(10);
	sub_wire2(143, 11)    <= sub_wire114(11);
	sub_wire2(143, 12)    <= sub_wire114(12);
	sub_wire2(143, 13)    <= sub_wire114(13);
	sub_wire2(143, 14)    <= sub_wire114(14);
	sub_wire2(143, 15)    <= sub_wire114(15);
	sub_wire2(143, 16)    <= sub_wire114(16);
	sub_wire2(143, 17)    <= sub_wire114(17);
	sub_wire2(143, 18)    <= sub_wire114(18);
	sub_wire2(143, 19)    <= sub_wire114(19);
	sub_wire2(143, 20)    <= sub_wire114(20);
	sub_wire2(143, 21)    <= sub_wire114(21);
	sub_wire2(143, 22)    <= sub_wire114(22);
	sub_wire2(143, 23)    <= sub_wire114(23);
	sub_wire2(143, 24)    <= sub_wire114(24);
	sub_wire2(143, 25)    <= sub_wire114(25);
	sub_wire2(143, 26)    <= sub_wire114(26);
	sub_wire2(143, 27)    <= sub_wire114(27);
	sub_wire2(143, 28)    <= sub_wire114(28);
	sub_wire2(143, 29)    <= sub_wire114(29);
	sub_wire2(143, 30)    <= sub_wire114(30);
	sub_wire2(143, 31)    <= sub_wire114(31);
	sub_wire2(143, 32)    <= sub_wire114(32);
	sub_wire2(143, 33)    <= sub_wire114(33);
	sub_wire2(143, 34)    <= sub_wire114(34);
	sub_wire2(143, 35)    <= sub_wire114(35);
	sub_wire2(143, 36)    <= sub_wire114(36);
	sub_wire2(143, 37)    <= sub_wire114(37);
	sub_wire2(143, 38)    <= sub_wire114(38);
	sub_wire2(143, 39)    <= sub_wire114(39);
	sub_wire2(142, 0)    <= sub_wire115(0);
	sub_wire2(142, 1)    <= sub_wire115(1);
	sub_wire2(142, 2)    <= sub_wire115(2);
	sub_wire2(142, 3)    <= sub_wire115(3);
	sub_wire2(142, 4)    <= sub_wire115(4);
	sub_wire2(142, 5)    <= sub_wire115(5);
	sub_wire2(142, 6)    <= sub_wire115(6);
	sub_wire2(142, 7)    <= sub_wire115(7);
	sub_wire2(142, 8)    <= sub_wire115(8);
	sub_wire2(142, 9)    <= sub_wire115(9);
	sub_wire2(142, 10)    <= sub_wire115(10);
	sub_wire2(142, 11)    <= sub_wire115(11);
	sub_wire2(142, 12)    <= sub_wire115(12);
	sub_wire2(142, 13)    <= sub_wire115(13);
	sub_wire2(142, 14)    <= sub_wire115(14);
	sub_wire2(142, 15)    <= sub_wire115(15);
	sub_wire2(142, 16)    <= sub_wire115(16);
	sub_wire2(142, 17)    <= sub_wire115(17);
	sub_wire2(142, 18)    <= sub_wire115(18);
	sub_wire2(142, 19)    <= sub_wire115(19);
	sub_wire2(142, 20)    <= sub_wire115(20);
	sub_wire2(142, 21)    <= sub_wire115(21);
	sub_wire2(142, 22)    <= sub_wire115(22);
	sub_wire2(142, 23)    <= sub_wire115(23);
	sub_wire2(142, 24)    <= sub_wire115(24);
	sub_wire2(142, 25)    <= sub_wire115(25);
	sub_wire2(142, 26)    <= sub_wire115(26);
	sub_wire2(142, 27)    <= sub_wire115(27);
	sub_wire2(142, 28)    <= sub_wire115(28);
	sub_wire2(142, 29)    <= sub_wire115(29);
	sub_wire2(142, 30)    <= sub_wire115(30);
	sub_wire2(142, 31)    <= sub_wire115(31);
	sub_wire2(142, 32)    <= sub_wire115(32);
	sub_wire2(142, 33)    <= sub_wire115(33);
	sub_wire2(142, 34)    <= sub_wire115(34);
	sub_wire2(142, 35)    <= sub_wire115(35);
	sub_wire2(142, 36)    <= sub_wire115(36);
	sub_wire2(142, 37)    <= sub_wire115(37);
	sub_wire2(142, 38)    <= sub_wire115(38);
	sub_wire2(142, 39)    <= sub_wire115(39);
	sub_wire2(141, 0)    <= sub_wire116(0);
	sub_wire2(141, 1)    <= sub_wire116(1);
	sub_wire2(141, 2)    <= sub_wire116(2);
	sub_wire2(141, 3)    <= sub_wire116(3);
	sub_wire2(141, 4)    <= sub_wire116(4);
	sub_wire2(141, 5)    <= sub_wire116(5);
	sub_wire2(141, 6)    <= sub_wire116(6);
	sub_wire2(141, 7)    <= sub_wire116(7);
	sub_wire2(141, 8)    <= sub_wire116(8);
	sub_wire2(141, 9)    <= sub_wire116(9);
	sub_wire2(141, 10)    <= sub_wire116(10);
	sub_wire2(141, 11)    <= sub_wire116(11);
	sub_wire2(141, 12)    <= sub_wire116(12);
	sub_wire2(141, 13)    <= sub_wire116(13);
	sub_wire2(141, 14)    <= sub_wire116(14);
	sub_wire2(141, 15)    <= sub_wire116(15);
	sub_wire2(141, 16)    <= sub_wire116(16);
	sub_wire2(141, 17)    <= sub_wire116(17);
	sub_wire2(141, 18)    <= sub_wire116(18);
	sub_wire2(141, 19)    <= sub_wire116(19);
	sub_wire2(141, 20)    <= sub_wire116(20);
	sub_wire2(141, 21)    <= sub_wire116(21);
	sub_wire2(141, 22)    <= sub_wire116(22);
	sub_wire2(141, 23)    <= sub_wire116(23);
	sub_wire2(141, 24)    <= sub_wire116(24);
	sub_wire2(141, 25)    <= sub_wire116(25);
	sub_wire2(141, 26)    <= sub_wire116(26);
	sub_wire2(141, 27)    <= sub_wire116(27);
	sub_wire2(141, 28)    <= sub_wire116(28);
	sub_wire2(141, 29)    <= sub_wire116(29);
	sub_wire2(141, 30)    <= sub_wire116(30);
	sub_wire2(141, 31)    <= sub_wire116(31);
	sub_wire2(141, 32)    <= sub_wire116(32);
	sub_wire2(141, 33)    <= sub_wire116(33);
	sub_wire2(141, 34)    <= sub_wire116(34);
	sub_wire2(141, 35)    <= sub_wire116(35);
	sub_wire2(141, 36)    <= sub_wire116(36);
	sub_wire2(141, 37)    <= sub_wire116(37);
	sub_wire2(141, 38)    <= sub_wire116(38);
	sub_wire2(141, 39)    <= sub_wire116(39);
	sub_wire2(140, 0)    <= sub_wire117(0);
	sub_wire2(140, 1)    <= sub_wire117(1);
	sub_wire2(140, 2)    <= sub_wire117(2);
	sub_wire2(140, 3)    <= sub_wire117(3);
	sub_wire2(140, 4)    <= sub_wire117(4);
	sub_wire2(140, 5)    <= sub_wire117(5);
	sub_wire2(140, 6)    <= sub_wire117(6);
	sub_wire2(140, 7)    <= sub_wire117(7);
	sub_wire2(140, 8)    <= sub_wire117(8);
	sub_wire2(140, 9)    <= sub_wire117(9);
	sub_wire2(140, 10)    <= sub_wire117(10);
	sub_wire2(140, 11)    <= sub_wire117(11);
	sub_wire2(140, 12)    <= sub_wire117(12);
	sub_wire2(140, 13)    <= sub_wire117(13);
	sub_wire2(140, 14)    <= sub_wire117(14);
	sub_wire2(140, 15)    <= sub_wire117(15);
	sub_wire2(140, 16)    <= sub_wire117(16);
	sub_wire2(140, 17)    <= sub_wire117(17);
	sub_wire2(140, 18)    <= sub_wire117(18);
	sub_wire2(140, 19)    <= sub_wire117(19);
	sub_wire2(140, 20)    <= sub_wire117(20);
	sub_wire2(140, 21)    <= sub_wire117(21);
	sub_wire2(140, 22)    <= sub_wire117(22);
	sub_wire2(140, 23)    <= sub_wire117(23);
	sub_wire2(140, 24)    <= sub_wire117(24);
	sub_wire2(140, 25)    <= sub_wire117(25);
	sub_wire2(140, 26)    <= sub_wire117(26);
	sub_wire2(140, 27)    <= sub_wire117(27);
	sub_wire2(140, 28)    <= sub_wire117(28);
	sub_wire2(140, 29)    <= sub_wire117(29);
	sub_wire2(140, 30)    <= sub_wire117(30);
	sub_wire2(140, 31)    <= sub_wire117(31);
	sub_wire2(140, 32)    <= sub_wire117(32);
	sub_wire2(140, 33)    <= sub_wire117(33);
	sub_wire2(140, 34)    <= sub_wire117(34);
	sub_wire2(140, 35)    <= sub_wire117(35);
	sub_wire2(140, 36)    <= sub_wire117(36);
	sub_wire2(140, 37)    <= sub_wire117(37);
	sub_wire2(140, 38)    <= sub_wire117(38);
	sub_wire2(140, 39)    <= sub_wire117(39);
	sub_wire2(139, 0)    <= sub_wire118(0);
	sub_wire2(139, 1)    <= sub_wire118(1);
	sub_wire2(139, 2)    <= sub_wire118(2);
	sub_wire2(139, 3)    <= sub_wire118(3);
	sub_wire2(139, 4)    <= sub_wire118(4);
	sub_wire2(139, 5)    <= sub_wire118(5);
	sub_wire2(139, 6)    <= sub_wire118(6);
	sub_wire2(139, 7)    <= sub_wire118(7);
	sub_wire2(139, 8)    <= sub_wire118(8);
	sub_wire2(139, 9)    <= sub_wire118(9);
	sub_wire2(139, 10)    <= sub_wire118(10);
	sub_wire2(139, 11)    <= sub_wire118(11);
	sub_wire2(139, 12)    <= sub_wire118(12);
	sub_wire2(139, 13)    <= sub_wire118(13);
	sub_wire2(139, 14)    <= sub_wire118(14);
	sub_wire2(139, 15)    <= sub_wire118(15);
	sub_wire2(139, 16)    <= sub_wire118(16);
	sub_wire2(139, 17)    <= sub_wire118(17);
	sub_wire2(139, 18)    <= sub_wire118(18);
	sub_wire2(139, 19)    <= sub_wire118(19);
	sub_wire2(139, 20)    <= sub_wire118(20);
	sub_wire2(139, 21)    <= sub_wire118(21);
	sub_wire2(139, 22)    <= sub_wire118(22);
	sub_wire2(139, 23)    <= sub_wire118(23);
	sub_wire2(139, 24)    <= sub_wire118(24);
	sub_wire2(139, 25)    <= sub_wire118(25);
	sub_wire2(139, 26)    <= sub_wire118(26);
	sub_wire2(139, 27)    <= sub_wire118(27);
	sub_wire2(139, 28)    <= sub_wire118(28);
	sub_wire2(139, 29)    <= sub_wire118(29);
	sub_wire2(139, 30)    <= sub_wire118(30);
	sub_wire2(139, 31)    <= sub_wire118(31);
	sub_wire2(139, 32)    <= sub_wire118(32);
	sub_wire2(139, 33)    <= sub_wire118(33);
	sub_wire2(139, 34)    <= sub_wire118(34);
	sub_wire2(139, 35)    <= sub_wire118(35);
	sub_wire2(139, 36)    <= sub_wire118(36);
	sub_wire2(139, 37)    <= sub_wire118(37);
	sub_wire2(139, 38)    <= sub_wire118(38);
	sub_wire2(139, 39)    <= sub_wire118(39);
	sub_wire2(138, 0)    <= sub_wire119(0);
	sub_wire2(138, 1)    <= sub_wire119(1);
	sub_wire2(138, 2)    <= sub_wire119(2);
	sub_wire2(138, 3)    <= sub_wire119(3);
	sub_wire2(138, 4)    <= sub_wire119(4);
	sub_wire2(138, 5)    <= sub_wire119(5);
	sub_wire2(138, 6)    <= sub_wire119(6);
	sub_wire2(138, 7)    <= sub_wire119(7);
	sub_wire2(138, 8)    <= sub_wire119(8);
	sub_wire2(138, 9)    <= sub_wire119(9);
	sub_wire2(138, 10)    <= sub_wire119(10);
	sub_wire2(138, 11)    <= sub_wire119(11);
	sub_wire2(138, 12)    <= sub_wire119(12);
	sub_wire2(138, 13)    <= sub_wire119(13);
	sub_wire2(138, 14)    <= sub_wire119(14);
	sub_wire2(138, 15)    <= sub_wire119(15);
	sub_wire2(138, 16)    <= sub_wire119(16);
	sub_wire2(138, 17)    <= sub_wire119(17);
	sub_wire2(138, 18)    <= sub_wire119(18);
	sub_wire2(138, 19)    <= sub_wire119(19);
	sub_wire2(138, 20)    <= sub_wire119(20);
	sub_wire2(138, 21)    <= sub_wire119(21);
	sub_wire2(138, 22)    <= sub_wire119(22);
	sub_wire2(138, 23)    <= sub_wire119(23);
	sub_wire2(138, 24)    <= sub_wire119(24);
	sub_wire2(138, 25)    <= sub_wire119(25);
	sub_wire2(138, 26)    <= sub_wire119(26);
	sub_wire2(138, 27)    <= sub_wire119(27);
	sub_wire2(138, 28)    <= sub_wire119(28);
	sub_wire2(138, 29)    <= sub_wire119(29);
	sub_wire2(138, 30)    <= sub_wire119(30);
	sub_wire2(138, 31)    <= sub_wire119(31);
	sub_wire2(138, 32)    <= sub_wire119(32);
	sub_wire2(138, 33)    <= sub_wire119(33);
	sub_wire2(138, 34)    <= sub_wire119(34);
	sub_wire2(138, 35)    <= sub_wire119(35);
	sub_wire2(138, 36)    <= sub_wire119(36);
	sub_wire2(138, 37)    <= sub_wire119(37);
	sub_wire2(138, 38)    <= sub_wire119(38);
	sub_wire2(138, 39)    <= sub_wire119(39);
	sub_wire2(137, 0)    <= sub_wire120(0);
	sub_wire2(137, 1)    <= sub_wire120(1);
	sub_wire2(137, 2)    <= sub_wire120(2);
	sub_wire2(137, 3)    <= sub_wire120(3);
	sub_wire2(137, 4)    <= sub_wire120(4);
	sub_wire2(137, 5)    <= sub_wire120(5);
	sub_wire2(137, 6)    <= sub_wire120(6);
	sub_wire2(137, 7)    <= sub_wire120(7);
	sub_wire2(137, 8)    <= sub_wire120(8);
	sub_wire2(137, 9)    <= sub_wire120(9);
	sub_wire2(137, 10)    <= sub_wire120(10);
	sub_wire2(137, 11)    <= sub_wire120(11);
	sub_wire2(137, 12)    <= sub_wire120(12);
	sub_wire2(137, 13)    <= sub_wire120(13);
	sub_wire2(137, 14)    <= sub_wire120(14);
	sub_wire2(137, 15)    <= sub_wire120(15);
	sub_wire2(137, 16)    <= sub_wire120(16);
	sub_wire2(137, 17)    <= sub_wire120(17);
	sub_wire2(137, 18)    <= sub_wire120(18);
	sub_wire2(137, 19)    <= sub_wire120(19);
	sub_wire2(137, 20)    <= sub_wire120(20);
	sub_wire2(137, 21)    <= sub_wire120(21);
	sub_wire2(137, 22)    <= sub_wire120(22);
	sub_wire2(137, 23)    <= sub_wire120(23);
	sub_wire2(137, 24)    <= sub_wire120(24);
	sub_wire2(137, 25)    <= sub_wire120(25);
	sub_wire2(137, 26)    <= sub_wire120(26);
	sub_wire2(137, 27)    <= sub_wire120(27);
	sub_wire2(137, 28)    <= sub_wire120(28);
	sub_wire2(137, 29)    <= sub_wire120(29);
	sub_wire2(137, 30)    <= sub_wire120(30);
	sub_wire2(137, 31)    <= sub_wire120(31);
	sub_wire2(137, 32)    <= sub_wire120(32);
	sub_wire2(137, 33)    <= sub_wire120(33);
	sub_wire2(137, 34)    <= sub_wire120(34);
	sub_wire2(137, 35)    <= sub_wire120(35);
	sub_wire2(137, 36)    <= sub_wire120(36);
	sub_wire2(137, 37)    <= sub_wire120(37);
	sub_wire2(137, 38)    <= sub_wire120(38);
	sub_wire2(137, 39)    <= sub_wire120(39);
	sub_wire2(136, 0)    <= sub_wire121(0);
	sub_wire2(136, 1)    <= sub_wire121(1);
	sub_wire2(136, 2)    <= sub_wire121(2);
	sub_wire2(136, 3)    <= sub_wire121(3);
	sub_wire2(136, 4)    <= sub_wire121(4);
	sub_wire2(136, 5)    <= sub_wire121(5);
	sub_wire2(136, 6)    <= sub_wire121(6);
	sub_wire2(136, 7)    <= sub_wire121(7);
	sub_wire2(136, 8)    <= sub_wire121(8);
	sub_wire2(136, 9)    <= sub_wire121(9);
	sub_wire2(136, 10)    <= sub_wire121(10);
	sub_wire2(136, 11)    <= sub_wire121(11);
	sub_wire2(136, 12)    <= sub_wire121(12);
	sub_wire2(136, 13)    <= sub_wire121(13);
	sub_wire2(136, 14)    <= sub_wire121(14);
	sub_wire2(136, 15)    <= sub_wire121(15);
	sub_wire2(136, 16)    <= sub_wire121(16);
	sub_wire2(136, 17)    <= sub_wire121(17);
	sub_wire2(136, 18)    <= sub_wire121(18);
	sub_wire2(136, 19)    <= sub_wire121(19);
	sub_wire2(136, 20)    <= sub_wire121(20);
	sub_wire2(136, 21)    <= sub_wire121(21);
	sub_wire2(136, 22)    <= sub_wire121(22);
	sub_wire2(136, 23)    <= sub_wire121(23);
	sub_wire2(136, 24)    <= sub_wire121(24);
	sub_wire2(136, 25)    <= sub_wire121(25);
	sub_wire2(136, 26)    <= sub_wire121(26);
	sub_wire2(136, 27)    <= sub_wire121(27);
	sub_wire2(136, 28)    <= sub_wire121(28);
	sub_wire2(136, 29)    <= sub_wire121(29);
	sub_wire2(136, 30)    <= sub_wire121(30);
	sub_wire2(136, 31)    <= sub_wire121(31);
	sub_wire2(136, 32)    <= sub_wire121(32);
	sub_wire2(136, 33)    <= sub_wire121(33);
	sub_wire2(136, 34)    <= sub_wire121(34);
	sub_wire2(136, 35)    <= sub_wire121(35);
	sub_wire2(136, 36)    <= sub_wire121(36);
	sub_wire2(136, 37)    <= sub_wire121(37);
	sub_wire2(136, 38)    <= sub_wire121(38);
	sub_wire2(136, 39)    <= sub_wire121(39);
	sub_wire2(135, 0)    <= sub_wire122(0);
	sub_wire2(135, 1)    <= sub_wire122(1);
	sub_wire2(135, 2)    <= sub_wire122(2);
	sub_wire2(135, 3)    <= sub_wire122(3);
	sub_wire2(135, 4)    <= sub_wire122(4);
	sub_wire2(135, 5)    <= sub_wire122(5);
	sub_wire2(135, 6)    <= sub_wire122(6);
	sub_wire2(135, 7)    <= sub_wire122(7);
	sub_wire2(135, 8)    <= sub_wire122(8);
	sub_wire2(135, 9)    <= sub_wire122(9);
	sub_wire2(135, 10)    <= sub_wire122(10);
	sub_wire2(135, 11)    <= sub_wire122(11);
	sub_wire2(135, 12)    <= sub_wire122(12);
	sub_wire2(135, 13)    <= sub_wire122(13);
	sub_wire2(135, 14)    <= sub_wire122(14);
	sub_wire2(135, 15)    <= sub_wire122(15);
	sub_wire2(135, 16)    <= sub_wire122(16);
	sub_wire2(135, 17)    <= sub_wire122(17);
	sub_wire2(135, 18)    <= sub_wire122(18);
	sub_wire2(135, 19)    <= sub_wire122(19);
	sub_wire2(135, 20)    <= sub_wire122(20);
	sub_wire2(135, 21)    <= sub_wire122(21);
	sub_wire2(135, 22)    <= sub_wire122(22);
	sub_wire2(135, 23)    <= sub_wire122(23);
	sub_wire2(135, 24)    <= sub_wire122(24);
	sub_wire2(135, 25)    <= sub_wire122(25);
	sub_wire2(135, 26)    <= sub_wire122(26);
	sub_wire2(135, 27)    <= sub_wire122(27);
	sub_wire2(135, 28)    <= sub_wire122(28);
	sub_wire2(135, 29)    <= sub_wire122(29);
	sub_wire2(135, 30)    <= sub_wire122(30);
	sub_wire2(135, 31)    <= sub_wire122(31);
	sub_wire2(135, 32)    <= sub_wire122(32);
	sub_wire2(135, 33)    <= sub_wire122(33);
	sub_wire2(135, 34)    <= sub_wire122(34);
	sub_wire2(135, 35)    <= sub_wire122(35);
	sub_wire2(135, 36)    <= sub_wire122(36);
	sub_wire2(135, 37)    <= sub_wire122(37);
	sub_wire2(135, 38)    <= sub_wire122(38);
	sub_wire2(135, 39)    <= sub_wire122(39);
	sub_wire2(134, 0)    <= sub_wire123(0);
	sub_wire2(134, 1)    <= sub_wire123(1);
	sub_wire2(134, 2)    <= sub_wire123(2);
	sub_wire2(134, 3)    <= sub_wire123(3);
	sub_wire2(134, 4)    <= sub_wire123(4);
	sub_wire2(134, 5)    <= sub_wire123(5);
	sub_wire2(134, 6)    <= sub_wire123(6);
	sub_wire2(134, 7)    <= sub_wire123(7);
	sub_wire2(134, 8)    <= sub_wire123(8);
	sub_wire2(134, 9)    <= sub_wire123(9);
	sub_wire2(134, 10)    <= sub_wire123(10);
	sub_wire2(134, 11)    <= sub_wire123(11);
	sub_wire2(134, 12)    <= sub_wire123(12);
	sub_wire2(134, 13)    <= sub_wire123(13);
	sub_wire2(134, 14)    <= sub_wire123(14);
	sub_wire2(134, 15)    <= sub_wire123(15);
	sub_wire2(134, 16)    <= sub_wire123(16);
	sub_wire2(134, 17)    <= sub_wire123(17);
	sub_wire2(134, 18)    <= sub_wire123(18);
	sub_wire2(134, 19)    <= sub_wire123(19);
	sub_wire2(134, 20)    <= sub_wire123(20);
	sub_wire2(134, 21)    <= sub_wire123(21);
	sub_wire2(134, 22)    <= sub_wire123(22);
	sub_wire2(134, 23)    <= sub_wire123(23);
	sub_wire2(134, 24)    <= sub_wire123(24);
	sub_wire2(134, 25)    <= sub_wire123(25);
	sub_wire2(134, 26)    <= sub_wire123(26);
	sub_wire2(134, 27)    <= sub_wire123(27);
	sub_wire2(134, 28)    <= sub_wire123(28);
	sub_wire2(134, 29)    <= sub_wire123(29);
	sub_wire2(134, 30)    <= sub_wire123(30);
	sub_wire2(134, 31)    <= sub_wire123(31);
	sub_wire2(134, 32)    <= sub_wire123(32);
	sub_wire2(134, 33)    <= sub_wire123(33);
	sub_wire2(134, 34)    <= sub_wire123(34);
	sub_wire2(134, 35)    <= sub_wire123(35);
	sub_wire2(134, 36)    <= sub_wire123(36);
	sub_wire2(134, 37)    <= sub_wire123(37);
	sub_wire2(134, 38)    <= sub_wire123(38);
	sub_wire2(134, 39)    <= sub_wire123(39);
	sub_wire2(133, 0)    <= sub_wire124(0);
	sub_wire2(133, 1)    <= sub_wire124(1);
	sub_wire2(133, 2)    <= sub_wire124(2);
	sub_wire2(133, 3)    <= sub_wire124(3);
	sub_wire2(133, 4)    <= sub_wire124(4);
	sub_wire2(133, 5)    <= sub_wire124(5);
	sub_wire2(133, 6)    <= sub_wire124(6);
	sub_wire2(133, 7)    <= sub_wire124(7);
	sub_wire2(133, 8)    <= sub_wire124(8);
	sub_wire2(133, 9)    <= sub_wire124(9);
	sub_wire2(133, 10)    <= sub_wire124(10);
	sub_wire2(133, 11)    <= sub_wire124(11);
	sub_wire2(133, 12)    <= sub_wire124(12);
	sub_wire2(133, 13)    <= sub_wire124(13);
	sub_wire2(133, 14)    <= sub_wire124(14);
	sub_wire2(133, 15)    <= sub_wire124(15);
	sub_wire2(133, 16)    <= sub_wire124(16);
	sub_wire2(133, 17)    <= sub_wire124(17);
	sub_wire2(133, 18)    <= sub_wire124(18);
	sub_wire2(133, 19)    <= sub_wire124(19);
	sub_wire2(133, 20)    <= sub_wire124(20);
	sub_wire2(133, 21)    <= sub_wire124(21);
	sub_wire2(133, 22)    <= sub_wire124(22);
	sub_wire2(133, 23)    <= sub_wire124(23);
	sub_wire2(133, 24)    <= sub_wire124(24);
	sub_wire2(133, 25)    <= sub_wire124(25);
	sub_wire2(133, 26)    <= sub_wire124(26);
	sub_wire2(133, 27)    <= sub_wire124(27);
	sub_wire2(133, 28)    <= sub_wire124(28);
	sub_wire2(133, 29)    <= sub_wire124(29);
	sub_wire2(133, 30)    <= sub_wire124(30);
	sub_wire2(133, 31)    <= sub_wire124(31);
	sub_wire2(133, 32)    <= sub_wire124(32);
	sub_wire2(133, 33)    <= sub_wire124(33);
	sub_wire2(133, 34)    <= sub_wire124(34);
	sub_wire2(133, 35)    <= sub_wire124(35);
	sub_wire2(133, 36)    <= sub_wire124(36);
	sub_wire2(133, 37)    <= sub_wire124(37);
	sub_wire2(133, 38)    <= sub_wire124(38);
	sub_wire2(133, 39)    <= sub_wire124(39);
	sub_wire2(132, 0)    <= sub_wire125(0);
	sub_wire2(132, 1)    <= sub_wire125(1);
	sub_wire2(132, 2)    <= sub_wire125(2);
	sub_wire2(132, 3)    <= sub_wire125(3);
	sub_wire2(132, 4)    <= sub_wire125(4);
	sub_wire2(132, 5)    <= sub_wire125(5);
	sub_wire2(132, 6)    <= sub_wire125(6);
	sub_wire2(132, 7)    <= sub_wire125(7);
	sub_wire2(132, 8)    <= sub_wire125(8);
	sub_wire2(132, 9)    <= sub_wire125(9);
	sub_wire2(132, 10)    <= sub_wire125(10);
	sub_wire2(132, 11)    <= sub_wire125(11);
	sub_wire2(132, 12)    <= sub_wire125(12);
	sub_wire2(132, 13)    <= sub_wire125(13);
	sub_wire2(132, 14)    <= sub_wire125(14);
	sub_wire2(132, 15)    <= sub_wire125(15);
	sub_wire2(132, 16)    <= sub_wire125(16);
	sub_wire2(132, 17)    <= sub_wire125(17);
	sub_wire2(132, 18)    <= sub_wire125(18);
	sub_wire2(132, 19)    <= sub_wire125(19);
	sub_wire2(132, 20)    <= sub_wire125(20);
	sub_wire2(132, 21)    <= sub_wire125(21);
	sub_wire2(132, 22)    <= sub_wire125(22);
	sub_wire2(132, 23)    <= sub_wire125(23);
	sub_wire2(132, 24)    <= sub_wire125(24);
	sub_wire2(132, 25)    <= sub_wire125(25);
	sub_wire2(132, 26)    <= sub_wire125(26);
	sub_wire2(132, 27)    <= sub_wire125(27);
	sub_wire2(132, 28)    <= sub_wire125(28);
	sub_wire2(132, 29)    <= sub_wire125(29);
	sub_wire2(132, 30)    <= sub_wire125(30);
	sub_wire2(132, 31)    <= sub_wire125(31);
	sub_wire2(132, 32)    <= sub_wire125(32);
	sub_wire2(132, 33)    <= sub_wire125(33);
	sub_wire2(132, 34)    <= sub_wire125(34);
	sub_wire2(132, 35)    <= sub_wire125(35);
	sub_wire2(132, 36)    <= sub_wire125(36);
	sub_wire2(132, 37)    <= sub_wire125(37);
	sub_wire2(132, 38)    <= sub_wire125(38);
	sub_wire2(132, 39)    <= sub_wire125(39);
	sub_wire2(131, 0)    <= sub_wire126(0);
	sub_wire2(131, 1)    <= sub_wire126(1);
	sub_wire2(131, 2)    <= sub_wire126(2);
	sub_wire2(131, 3)    <= sub_wire126(3);
	sub_wire2(131, 4)    <= sub_wire126(4);
	sub_wire2(131, 5)    <= sub_wire126(5);
	sub_wire2(131, 6)    <= sub_wire126(6);
	sub_wire2(131, 7)    <= sub_wire126(7);
	sub_wire2(131, 8)    <= sub_wire126(8);
	sub_wire2(131, 9)    <= sub_wire126(9);
	sub_wire2(131, 10)    <= sub_wire126(10);
	sub_wire2(131, 11)    <= sub_wire126(11);
	sub_wire2(131, 12)    <= sub_wire126(12);
	sub_wire2(131, 13)    <= sub_wire126(13);
	sub_wire2(131, 14)    <= sub_wire126(14);
	sub_wire2(131, 15)    <= sub_wire126(15);
	sub_wire2(131, 16)    <= sub_wire126(16);
	sub_wire2(131, 17)    <= sub_wire126(17);
	sub_wire2(131, 18)    <= sub_wire126(18);
	sub_wire2(131, 19)    <= sub_wire126(19);
	sub_wire2(131, 20)    <= sub_wire126(20);
	sub_wire2(131, 21)    <= sub_wire126(21);
	sub_wire2(131, 22)    <= sub_wire126(22);
	sub_wire2(131, 23)    <= sub_wire126(23);
	sub_wire2(131, 24)    <= sub_wire126(24);
	sub_wire2(131, 25)    <= sub_wire126(25);
	sub_wire2(131, 26)    <= sub_wire126(26);
	sub_wire2(131, 27)    <= sub_wire126(27);
	sub_wire2(131, 28)    <= sub_wire126(28);
	sub_wire2(131, 29)    <= sub_wire126(29);
	sub_wire2(131, 30)    <= sub_wire126(30);
	sub_wire2(131, 31)    <= sub_wire126(31);
	sub_wire2(131, 32)    <= sub_wire126(32);
	sub_wire2(131, 33)    <= sub_wire126(33);
	sub_wire2(131, 34)    <= sub_wire126(34);
	sub_wire2(131, 35)    <= sub_wire126(35);
	sub_wire2(131, 36)    <= sub_wire126(36);
	sub_wire2(131, 37)    <= sub_wire126(37);
	sub_wire2(131, 38)    <= sub_wire126(38);
	sub_wire2(131, 39)    <= sub_wire126(39);
	sub_wire2(130, 0)    <= sub_wire127(0);
	sub_wire2(130, 1)    <= sub_wire127(1);
	sub_wire2(130, 2)    <= sub_wire127(2);
	sub_wire2(130, 3)    <= sub_wire127(3);
	sub_wire2(130, 4)    <= sub_wire127(4);
	sub_wire2(130, 5)    <= sub_wire127(5);
	sub_wire2(130, 6)    <= sub_wire127(6);
	sub_wire2(130, 7)    <= sub_wire127(7);
	sub_wire2(130, 8)    <= sub_wire127(8);
	sub_wire2(130, 9)    <= sub_wire127(9);
	sub_wire2(130, 10)    <= sub_wire127(10);
	sub_wire2(130, 11)    <= sub_wire127(11);
	sub_wire2(130, 12)    <= sub_wire127(12);
	sub_wire2(130, 13)    <= sub_wire127(13);
	sub_wire2(130, 14)    <= sub_wire127(14);
	sub_wire2(130, 15)    <= sub_wire127(15);
	sub_wire2(130, 16)    <= sub_wire127(16);
	sub_wire2(130, 17)    <= sub_wire127(17);
	sub_wire2(130, 18)    <= sub_wire127(18);
	sub_wire2(130, 19)    <= sub_wire127(19);
	sub_wire2(130, 20)    <= sub_wire127(20);
	sub_wire2(130, 21)    <= sub_wire127(21);
	sub_wire2(130, 22)    <= sub_wire127(22);
	sub_wire2(130, 23)    <= sub_wire127(23);
	sub_wire2(130, 24)    <= sub_wire127(24);
	sub_wire2(130, 25)    <= sub_wire127(25);
	sub_wire2(130, 26)    <= sub_wire127(26);
	sub_wire2(130, 27)    <= sub_wire127(27);
	sub_wire2(130, 28)    <= sub_wire127(28);
	sub_wire2(130, 29)    <= sub_wire127(29);
	sub_wire2(130, 30)    <= sub_wire127(30);
	sub_wire2(130, 31)    <= sub_wire127(31);
	sub_wire2(130, 32)    <= sub_wire127(32);
	sub_wire2(130, 33)    <= sub_wire127(33);
	sub_wire2(130, 34)    <= sub_wire127(34);
	sub_wire2(130, 35)    <= sub_wire127(35);
	sub_wire2(130, 36)    <= sub_wire127(36);
	sub_wire2(130, 37)    <= sub_wire127(37);
	sub_wire2(130, 38)    <= sub_wire127(38);
	sub_wire2(130, 39)    <= sub_wire127(39);
	sub_wire2(129, 0)    <= sub_wire128(0);
	sub_wire2(129, 1)    <= sub_wire128(1);
	sub_wire2(129, 2)    <= sub_wire128(2);
	sub_wire2(129, 3)    <= sub_wire128(3);
	sub_wire2(129, 4)    <= sub_wire128(4);
	sub_wire2(129, 5)    <= sub_wire128(5);
	sub_wire2(129, 6)    <= sub_wire128(6);
	sub_wire2(129, 7)    <= sub_wire128(7);
	sub_wire2(129, 8)    <= sub_wire128(8);
	sub_wire2(129, 9)    <= sub_wire128(9);
	sub_wire2(129, 10)    <= sub_wire128(10);
	sub_wire2(129, 11)    <= sub_wire128(11);
	sub_wire2(129, 12)    <= sub_wire128(12);
	sub_wire2(129, 13)    <= sub_wire128(13);
	sub_wire2(129, 14)    <= sub_wire128(14);
	sub_wire2(129, 15)    <= sub_wire128(15);
	sub_wire2(129, 16)    <= sub_wire128(16);
	sub_wire2(129, 17)    <= sub_wire128(17);
	sub_wire2(129, 18)    <= sub_wire128(18);
	sub_wire2(129, 19)    <= sub_wire128(19);
	sub_wire2(129, 20)    <= sub_wire128(20);
	sub_wire2(129, 21)    <= sub_wire128(21);
	sub_wire2(129, 22)    <= sub_wire128(22);
	sub_wire2(129, 23)    <= sub_wire128(23);
	sub_wire2(129, 24)    <= sub_wire128(24);
	sub_wire2(129, 25)    <= sub_wire128(25);
	sub_wire2(129, 26)    <= sub_wire128(26);
	sub_wire2(129, 27)    <= sub_wire128(27);
	sub_wire2(129, 28)    <= sub_wire128(28);
	sub_wire2(129, 29)    <= sub_wire128(29);
	sub_wire2(129, 30)    <= sub_wire128(30);
	sub_wire2(129, 31)    <= sub_wire128(31);
	sub_wire2(129, 32)    <= sub_wire128(32);
	sub_wire2(129, 33)    <= sub_wire128(33);
	sub_wire2(129, 34)    <= sub_wire128(34);
	sub_wire2(129, 35)    <= sub_wire128(35);
	sub_wire2(129, 36)    <= sub_wire128(36);
	sub_wire2(129, 37)    <= sub_wire128(37);
	sub_wire2(129, 38)    <= sub_wire128(38);
	sub_wire2(129, 39)    <= sub_wire128(39);
	sub_wire2(128, 0)    <= sub_wire129(0);
	sub_wire2(128, 1)    <= sub_wire129(1);
	sub_wire2(128, 2)    <= sub_wire129(2);
	sub_wire2(128, 3)    <= sub_wire129(3);
	sub_wire2(128, 4)    <= sub_wire129(4);
	sub_wire2(128, 5)    <= sub_wire129(5);
	sub_wire2(128, 6)    <= sub_wire129(6);
	sub_wire2(128, 7)    <= sub_wire129(7);
	sub_wire2(128, 8)    <= sub_wire129(8);
	sub_wire2(128, 9)    <= sub_wire129(9);
	sub_wire2(128, 10)    <= sub_wire129(10);
	sub_wire2(128, 11)    <= sub_wire129(11);
	sub_wire2(128, 12)    <= sub_wire129(12);
	sub_wire2(128, 13)    <= sub_wire129(13);
	sub_wire2(128, 14)    <= sub_wire129(14);
	sub_wire2(128, 15)    <= sub_wire129(15);
	sub_wire2(128, 16)    <= sub_wire129(16);
	sub_wire2(128, 17)    <= sub_wire129(17);
	sub_wire2(128, 18)    <= sub_wire129(18);
	sub_wire2(128, 19)    <= sub_wire129(19);
	sub_wire2(128, 20)    <= sub_wire129(20);
	sub_wire2(128, 21)    <= sub_wire129(21);
	sub_wire2(128, 22)    <= sub_wire129(22);
	sub_wire2(128, 23)    <= sub_wire129(23);
	sub_wire2(128, 24)    <= sub_wire129(24);
	sub_wire2(128, 25)    <= sub_wire129(25);
	sub_wire2(128, 26)    <= sub_wire129(26);
	sub_wire2(128, 27)    <= sub_wire129(27);
	sub_wire2(128, 28)    <= sub_wire129(28);
	sub_wire2(128, 29)    <= sub_wire129(29);
	sub_wire2(128, 30)    <= sub_wire129(30);
	sub_wire2(128, 31)    <= sub_wire129(31);
	sub_wire2(128, 32)    <= sub_wire129(32);
	sub_wire2(128, 33)    <= sub_wire129(33);
	sub_wire2(128, 34)    <= sub_wire129(34);
	sub_wire2(128, 35)    <= sub_wire129(35);
	sub_wire2(128, 36)    <= sub_wire129(36);
	sub_wire2(128, 37)    <= sub_wire129(37);
	sub_wire2(128, 38)    <= sub_wire129(38);
	sub_wire2(128, 39)    <= sub_wire129(39);
	sub_wire2(127, 0)    <= sub_wire130(0);
	sub_wire2(127, 1)    <= sub_wire130(1);
	sub_wire2(127, 2)    <= sub_wire130(2);
	sub_wire2(127, 3)    <= sub_wire130(3);
	sub_wire2(127, 4)    <= sub_wire130(4);
	sub_wire2(127, 5)    <= sub_wire130(5);
	sub_wire2(127, 6)    <= sub_wire130(6);
	sub_wire2(127, 7)    <= sub_wire130(7);
	sub_wire2(127, 8)    <= sub_wire130(8);
	sub_wire2(127, 9)    <= sub_wire130(9);
	sub_wire2(127, 10)    <= sub_wire130(10);
	sub_wire2(127, 11)    <= sub_wire130(11);
	sub_wire2(127, 12)    <= sub_wire130(12);
	sub_wire2(127, 13)    <= sub_wire130(13);
	sub_wire2(127, 14)    <= sub_wire130(14);
	sub_wire2(127, 15)    <= sub_wire130(15);
	sub_wire2(127, 16)    <= sub_wire130(16);
	sub_wire2(127, 17)    <= sub_wire130(17);
	sub_wire2(127, 18)    <= sub_wire130(18);
	sub_wire2(127, 19)    <= sub_wire130(19);
	sub_wire2(127, 20)    <= sub_wire130(20);
	sub_wire2(127, 21)    <= sub_wire130(21);
	sub_wire2(127, 22)    <= sub_wire130(22);
	sub_wire2(127, 23)    <= sub_wire130(23);
	sub_wire2(127, 24)    <= sub_wire130(24);
	sub_wire2(127, 25)    <= sub_wire130(25);
	sub_wire2(127, 26)    <= sub_wire130(26);
	sub_wire2(127, 27)    <= sub_wire130(27);
	sub_wire2(127, 28)    <= sub_wire130(28);
	sub_wire2(127, 29)    <= sub_wire130(29);
	sub_wire2(127, 30)    <= sub_wire130(30);
	sub_wire2(127, 31)    <= sub_wire130(31);
	sub_wire2(127, 32)    <= sub_wire130(32);
	sub_wire2(127, 33)    <= sub_wire130(33);
	sub_wire2(127, 34)    <= sub_wire130(34);
	sub_wire2(127, 35)    <= sub_wire130(35);
	sub_wire2(127, 36)    <= sub_wire130(36);
	sub_wire2(127, 37)    <= sub_wire130(37);
	sub_wire2(127, 38)    <= sub_wire130(38);
	sub_wire2(127, 39)    <= sub_wire130(39);
	sub_wire2(126, 0)    <= sub_wire131(0);
	sub_wire2(126, 1)    <= sub_wire131(1);
	sub_wire2(126, 2)    <= sub_wire131(2);
	sub_wire2(126, 3)    <= sub_wire131(3);
	sub_wire2(126, 4)    <= sub_wire131(4);
	sub_wire2(126, 5)    <= sub_wire131(5);
	sub_wire2(126, 6)    <= sub_wire131(6);
	sub_wire2(126, 7)    <= sub_wire131(7);
	sub_wire2(126, 8)    <= sub_wire131(8);
	sub_wire2(126, 9)    <= sub_wire131(9);
	sub_wire2(126, 10)    <= sub_wire131(10);
	sub_wire2(126, 11)    <= sub_wire131(11);
	sub_wire2(126, 12)    <= sub_wire131(12);
	sub_wire2(126, 13)    <= sub_wire131(13);
	sub_wire2(126, 14)    <= sub_wire131(14);
	sub_wire2(126, 15)    <= sub_wire131(15);
	sub_wire2(126, 16)    <= sub_wire131(16);
	sub_wire2(126, 17)    <= sub_wire131(17);
	sub_wire2(126, 18)    <= sub_wire131(18);
	sub_wire2(126, 19)    <= sub_wire131(19);
	sub_wire2(126, 20)    <= sub_wire131(20);
	sub_wire2(126, 21)    <= sub_wire131(21);
	sub_wire2(126, 22)    <= sub_wire131(22);
	sub_wire2(126, 23)    <= sub_wire131(23);
	sub_wire2(126, 24)    <= sub_wire131(24);
	sub_wire2(126, 25)    <= sub_wire131(25);
	sub_wire2(126, 26)    <= sub_wire131(26);
	sub_wire2(126, 27)    <= sub_wire131(27);
	sub_wire2(126, 28)    <= sub_wire131(28);
	sub_wire2(126, 29)    <= sub_wire131(29);
	sub_wire2(126, 30)    <= sub_wire131(30);
	sub_wire2(126, 31)    <= sub_wire131(31);
	sub_wire2(126, 32)    <= sub_wire131(32);
	sub_wire2(126, 33)    <= sub_wire131(33);
	sub_wire2(126, 34)    <= sub_wire131(34);
	sub_wire2(126, 35)    <= sub_wire131(35);
	sub_wire2(126, 36)    <= sub_wire131(36);
	sub_wire2(126, 37)    <= sub_wire131(37);
	sub_wire2(126, 38)    <= sub_wire131(38);
	sub_wire2(126, 39)    <= sub_wire131(39);
	sub_wire2(125, 0)    <= sub_wire132(0);
	sub_wire2(125, 1)    <= sub_wire132(1);
	sub_wire2(125, 2)    <= sub_wire132(2);
	sub_wire2(125, 3)    <= sub_wire132(3);
	sub_wire2(125, 4)    <= sub_wire132(4);
	sub_wire2(125, 5)    <= sub_wire132(5);
	sub_wire2(125, 6)    <= sub_wire132(6);
	sub_wire2(125, 7)    <= sub_wire132(7);
	sub_wire2(125, 8)    <= sub_wire132(8);
	sub_wire2(125, 9)    <= sub_wire132(9);
	sub_wire2(125, 10)    <= sub_wire132(10);
	sub_wire2(125, 11)    <= sub_wire132(11);
	sub_wire2(125, 12)    <= sub_wire132(12);
	sub_wire2(125, 13)    <= sub_wire132(13);
	sub_wire2(125, 14)    <= sub_wire132(14);
	sub_wire2(125, 15)    <= sub_wire132(15);
	sub_wire2(125, 16)    <= sub_wire132(16);
	sub_wire2(125, 17)    <= sub_wire132(17);
	sub_wire2(125, 18)    <= sub_wire132(18);
	sub_wire2(125, 19)    <= sub_wire132(19);
	sub_wire2(125, 20)    <= sub_wire132(20);
	sub_wire2(125, 21)    <= sub_wire132(21);
	sub_wire2(125, 22)    <= sub_wire132(22);
	sub_wire2(125, 23)    <= sub_wire132(23);
	sub_wire2(125, 24)    <= sub_wire132(24);
	sub_wire2(125, 25)    <= sub_wire132(25);
	sub_wire2(125, 26)    <= sub_wire132(26);
	sub_wire2(125, 27)    <= sub_wire132(27);
	sub_wire2(125, 28)    <= sub_wire132(28);
	sub_wire2(125, 29)    <= sub_wire132(29);
	sub_wire2(125, 30)    <= sub_wire132(30);
	sub_wire2(125, 31)    <= sub_wire132(31);
	sub_wire2(125, 32)    <= sub_wire132(32);
	sub_wire2(125, 33)    <= sub_wire132(33);
	sub_wire2(125, 34)    <= sub_wire132(34);
	sub_wire2(125, 35)    <= sub_wire132(35);
	sub_wire2(125, 36)    <= sub_wire132(36);
	sub_wire2(125, 37)    <= sub_wire132(37);
	sub_wire2(125, 38)    <= sub_wire132(38);
	sub_wire2(125, 39)    <= sub_wire132(39);
	sub_wire2(124, 0)    <= sub_wire133(0);
	sub_wire2(124, 1)    <= sub_wire133(1);
	sub_wire2(124, 2)    <= sub_wire133(2);
	sub_wire2(124, 3)    <= sub_wire133(3);
	sub_wire2(124, 4)    <= sub_wire133(4);
	sub_wire2(124, 5)    <= sub_wire133(5);
	sub_wire2(124, 6)    <= sub_wire133(6);
	sub_wire2(124, 7)    <= sub_wire133(7);
	sub_wire2(124, 8)    <= sub_wire133(8);
	sub_wire2(124, 9)    <= sub_wire133(9);
	sub_wire2(124, 10)    <= sub_wire133(10);
	sub_wire2(124, 11)    <= sub_wire133(11);
	sub_wire2(124, 12)    <= sub_wire133(12);
	sub_wire2(124, 13)    <= sub_wire133(13);
	sub_wire2(124, 14)    <= sub_wire133(14);
	sub_wire2(124, 15)    <= sub_wire133(15);
	sub_wire2(124, 16)    <= sub_wire133(16);
	sub_wire2(124, 17)    <= sub_wire133(17);
	sub_wire2(124, 18)    <= sub_wire133(18);
	sub_wire2(124, 19)    <= sub_wire133(19);
	sub_wire2(124, 20)    <= sub_wire133(20);
	sub_wire2(124, 21)    <= sub_wire133(21);
	sub_wire2(124, 22)    <= sub_wire133(22);
	sub_wire2(124, 23)    <= sub_wire133(23);
	sub_wire2(124, 24)    <= sub_wire133(24);
	sub_wire2(124, 25)    <= sub_wire133(25);
	sub_wire2(124, 26)    <= sub_wire133(26);
	sub_wire2(124, 27)    <= sub_wire133(27);
	sub_wire2(124, 28)    <= sub_wire133(28);
	sub_wire2(124, 29)    <= sub_wire133(29);
	sub_wire2(124, 30)    <= sub_wire133(30);
	sub_wire2(124, 31)    <= sub_wire133(31);
	sub_wire2(124, 32)    <= sub_wire133(32);
	sub_wire2(124, 33)    <= sub_wire133(33);
	sub_wire2(124, 34)    <= sub_wire133(34);
	sub_wire2(124, 35)    <= sub_wire133(35);
	sub_wire2(124, 36)    <= sub_wire133(36);
	sub_wire2(124, 37)    <= sub_wire133(37);
	sub_wire2(124, 38)    <= sub_wire133(38);
	sub_wire2(124, 39)    <= sub_wire133(39);
	sub_wire2(123, 0)    <= sub_wire134(0);
	sub_wire2(123, 1)    <= sub_wire134(1);
	sub_wire2(123, 2)    <= sub_wire134(2);
	sub_wire2(123, 3)    <= sub_wire134(3);
	sub_wire2(123, 4)    <= sub_wire134(4);
	sub_wire2(123, 5)    <= sub_wire134(5);
	sub_wire2(123, 6)    <= sub_wire134(6);
	sub_wire2(123, 7)    <= sub_wire134(7);
	sub_wire2(123, 8)    <= sub_wire134(8);
	sub_wire2(123, 9)    <= sub_wire134(9);
	sub_wire2(123, 10)    <= sub_wire134(10);
	sub_wire2(123, 11)    <= sub_wire134(11);
	sub_wire2(123, 12)    <= sub_wire134(12);
	sub_wire2(123, 13)    <= sub_wire134(13);
	sub_wire2(123, 14)    <= sub_wire134(14);
	sub_wire2(123, 15)    <= sub_wire134(15);
	sub_wire2(123, 16)    <= sub_wire134(16);
	sub_wire2(123, 17)    <= sub_wire134(17);
	sub_wire2(123, 18)    <= sub_wire134(18);
	sub_wire2(123, 19)    <= sub_wire134(19);
	sub_wire2(123, 20)    <= sub_wire134(20);
	sub_wire2(123, 21)    <= sub_wire134(21);
	sub_wire2(123, 22)    <= sub_wire134(22);
	sub_wire2(123, 23)    <= sub_wire134(23);
	sub_wire2(123, 24)    <= sub_wire134(24);
	sub_wire2(123, 25)    <= sub_wire134(25);
	sub_wire2(123, 26)    <= sub_wire134(26);
	sub_wire2(123, 27)    <= sub_wire134(27);
	sub_wire2(123, 28)    <= sub_wire134(28);
	sub_wire2(123, 29)    <= sub_wire134(29);
	sub_wire2(123, 30)    <= sub_wire134(30);
	sub_wire2(123, 31)    <= sub_wire134(31);
	sub_wire2(123, 32)    <= sub_wire134(32);
	sub_wire2(123, 33)    <= sub_wire134(33);
	sub_wire2(123, 34)    <= sub_wire134(34);
	sub_wire2(123, 35)    <= sub_wire134(35);
	sub_wire2(123, 36)    <= sub_wire134(36);
	sub_wire2(123, 37)    <= sub_wire134(37);
	sub_wire2(123, 38)    <= sub_wire134(38);
	sub_wire2(123, 39)    <= sub_wire134(39);
	sub_wire2(122, 0)    <= sub_wire135(0);
	sub_wire2(122, 1)    <= sub_wire135(1);
	sub_wire2(122, 2)    <= sub_wire135(2);
	sub_wire2(122, 3)    <= sub_wire135(3);
	sub_wire2(122, 4)    <= sub_wire135(4);
	sub_wire2(122, 5)    <= sub_wire135(5);
	sub_wire2(122, 6)    <= sub_wire135(6);
	sub_wire2(122, 7)    <= sub_wire135(7);
	sub_wire2(122, 8)    <= sub_wire135(8);
	sub_wire2(122, 9)    <= sub_wire135(9);
	sub_wire2(122, 10)    <= sub_wire135(10);
	sub_wire2(122, 11)    <= sub_wire135(11);
	sub_wire2(122, 12)    <= sub_wire135(12);
	sub_wire2(122, 13)    <= sub_wire135(13);
	sub_wire2(122, 14)    <= sub_wire135(14);
	sub_wire2(122, 15)    <= sub_wire135(15);
	sub_wire2(122, 16)    <= sub_wire135(16);
	sub_wire2(122, 17)    <= sub_wire135(17);
	sub_wire2(122, 18)    <= sub_wire135(18);
	sub_wire2(122, 19)    <= sub_wire135(19);
	sub_wire2(122, 20)    <= sub_wire135(20);
	sub_wire2(122, 21)    <= sub_wire135(21);
	sub_wire2(122, 22)    <= sub_wire135(22);
	sub_wire2(122, 23)    <= sub_wire135(23);
	sub_wire2(122, 24)    <= sub_wire135(24);
	sub_wire2(122, 25)    <= sub_wire135(25);
	sub_wire2(122, 26)    <= sub_wire135(26);
	sub_wire2(122, 27)    <= sub_wire135(27);
	sub_wire2(122, 28)    <= sub_wire135(28);
	sub_wire2(122, 29)    <= sub_wire135(29);
	sub_wire2(122, 30)    <= sub_wire135(30);
	sub_wire2(122, 31)    <= sub_wire135(31);
	sub_wire2(122, 32)    <= sub_wire135(32);
	sub_wire2(122, 33)    <= sub_wire135(33);
	sub_wire2(122, 34)    <= sub_wire135(34);
	sub_wire2(122, 35)    <= sub_wire135(35);
	sub_wire2(122, 36)    <= sub_wire135(36);
	sub_wire2(122, 37)    <= sub_wire135(37);
	sub_wire2(122, 38)    <= sub_wire135(38);
	sub_wire2(122, 39)    <= sub_wire135(39);
	sub_wire2(121, 0)    <= sub_wire136(0);
	sub_wire2(121, 1)    <= sub_wire136(1);
	sub_wire2(121, 2)    <= sub_wire136(2);
	sub_wire2(121, 3)    <= sub_wire136(3);
	sub_wire2(121, 4)    <= sub_wire136(4);
	sub_wire2(121, 5)    <= sub_wire136(5);
	sub_wire2(121, 6)    <= sub_wire136(6);
	sub_wire2(121, 7)    <= sub_wire136(7);
	sub_wire2(121, 8)    <= sub_wire136(8);
	sub_wire2(121, 9)    <= sub_wire136(9);
	sub_wire2(121, 10)    <= sub_wire136(10);
	sub_wire2(121, 11)    <= sub_wire136(11);
	sub_wire2(121, 12)    <= sub_wire136(12);
	sub_wire2(121, 13)    <= sub_wire136(13);
	sub_wire2(121, 14)    <= sub_wire136(14);
	sub_wire2(121, 15)    <= sub_wire136(15);
	sub_wire2(121, 16)    <= sub_wire136(16);
	sub_wire2(121, 17)    <= sub_wire136(17);
	sub_wire2(121, 18)    <= sub_wire136(18);
	sub_wire2(121, 19)    <= sub_wire136(19);
	sub_wire2(121, 20)    <= sub_wire136(20);
	sub_wire2(121, 21)    <= sub_wire136(21);
	sub_wire2(121, 22)    <= sub_wire136(22);
	sub_wire2(121, 23)    <= sub_wire136(23);
	sub_wire2(121, 24)    <= sub_wire136(24);
	sub_wire2(121, 25)    <= sub_wire136(25);
	sub_wire2(121, 26)    <= sub_wire136(26);
	sub_wire2(121, 27)    <= sub_wire136(27);
	sub_wire2(121, 28)    <= sub_wire136(28);
	sub_wire2(121, 29)    <= sub_wire136(29);
	sub_wire2(121, 30)    <= sub_wire136(30);
	sub_wire2(121, 31)    <= sub_wire136(31);
	sub_wire2(121, 32)    <= sub_wire136(32);
	sub_wire2(121, 33)    <= sub_wire136(33);
	sub_wire2(121, 34)    <= sub_wire136(34);
	sub_wire2(121, 35)    <= sub_wire136(35);
	sub_wire2(121, 36)    <= sub_wire136(36);
	sub_wire2(121, 37)    <= sub_wire136(37);
	sub_wire2(121, 38)    <= sub_wire136(38);
	sub_wire2(121, 39)    <= sub_wire136(39);
	sub_wire2(120, 0)    <= sub_wire137(0);
	sub_wire2(120, 1)    <= sub_wire137(1);
	sub_wire2(120, 2)    <= sub_wire137(2);
	sub_wire2(120, 3)    <= sub_wire137(3);
	sub_wire2(120, 4)    <= sub_wire137(4);
	sub_wire2(120, 5)    <= sub_wire137(5);
	sub_wire2(120, 6)    <= sub_wire137(6);
	sub_wire2(120, 7)    <= sub_wire137(7);
	sub_wire2(120, 8)    <= sub_wire137(8);
	sub_wire2(120, 9)    <= sub_wire137(9);
	sub_wire2(120, 10)    <= sub_wire137(10);
	sub_wire2(120, 11)    <= sub_wire137(11);
	sub_wire2(120, 12)    <= sub_wire137(12);
	sub_wire2(120, 13)    <= sub_wire137(13);
	sub_wire2(120, 14)    <= sub_wire137(14);
	sub_wire2(120, 15)    <= sub_wire137(15);
	sub_wire2(120, 16)    <= sub_wire137(16);
	sub_wire2(120, 17)    <= sub_wire137(17);
	sub_wire2(120, 18)    <= sub_wire137(18);
	sub_wire2(120, 19)    <= sub_wire137(19);
	sub_wire2(120, 20)    <= sub_wire137(20);
	sub_wire2(120, 21)    <= sub_wire137(21);
	sub_wire2(120, 22)    <= sub_wire137(22);
	sub_wire2(120, 23)    <= sub_wire137(23);
	sub_wire2(120, 24)    <= sub_wire137(24);
	sub_wire2(120, 25)    <= sub_wire137(25);
	sub_wire2(120, 26)    <= sub_wire137(26);
	sub_wire2(120, 27)    <= sub_wire137(27);
	sub_wire2(120, 28)    <= sub_wire137(28);
	sub_wire2(120, 29)    <= sub_wire137(29);
	sub_wire2(120, 30)    <= sub_wire137(30);
	sub_wire2(120, 31)    <= sub_wire137(31);
	sub_wire2(120, 32)    <= sub_wire137(32);
	sub_wire2(120, 33)    <= sub_wire137(33);
	sub_wire2(120, 34)    <= sub_wire137(34);
	sub_wire2(120, 35)    <= sub_wire137(35);
	sub_wire2(120, 36)    <= sub_wire137(36);
	sub_wire2(120, 37)    <= sub_wire137(37);
	sub_wire2(120, 38)    <= sub_wire137(38);
	sub_wire2(120, 39)    <= sub_wire137(39);
	sub_wire2(119, 0)    <= sub_wire138(0);
	sub_wire2(119, 1)    <= sub_wire138(1);
	sub_wire2(119, 2)    <= sub_wire138(2);
	sub_wire2(119, 3)    <= sub_wire138(3);
	sub_wire2(119, 4)    <= sub_wire138(4);
	sub_wire2(119, 5)    <= sub_wire138(5);
	sub_wire2(119, 6)    <= sub_wire138(6);
	sub_wire2(119, 7)    <= sub_wire138(7);
	sub_wire2(119, 8)    <= sub_wire138(8);
	sub_wire2(119, 9)    <= sub_wire138(9);
	sub_wire2(119, 10)    <= sub_wire138(10);
	sub_wire2(119, 11)    <= sub_wire138(11);
	sub_wire2(119, 12)    <= sub_wire138(12);
	sub_wire2(119, 13)    <= sub_wire138(13);
	sub_wire2(119, 14)    <= sub_wire138(14);
	sub_wire2(119, 15)    <= sub_wire138(15);
	sub_wire2(119, 16)    <= sub_wire138(16);
	sub_wire2(119, 17)    <= sub_wire138(17);
	sub_wire2(119, 18)    <= sub_wire138(18);
	sub_wire2(119, 19)    <= sub_wire138(19);
	sub_wire2(119, 20)    <= sub_wire138(20);
	sub_wire2(119, 21)    <= sub_wire138(21);
	sub_wire2(119, 22)    <= sub_wire138(22);
	sub_wire2(119, 23)    <= sub_wire138(23);
	sub_wire2(119, 24)    <= sub_wire138(24);
	sub_wire2(119, 25)    <= sub_wire138(25);
	sub_wire2(119, 26)    <= sub_wire138(26);
	sub_wire2(119, 27)    <= sub_wire138(27);
	sub_wire2(119, 28)    <= sub_wire138(28);
	sub_wire2(119, 29)    <= sub_wire138(29);
	sub_wire2(119, 30)    <= sub_wire138(30);
	sub_wire2(119, 31)    <= sub_wire138(31);
	sub_wire2(119, 32)    <= sub_wire138(32);
	sub_wire2(119, 33)    <= sub_wire138(33);
	sub_wire2(119, 34)    <= sub_wire138(34);
	sub_wire2(119, 35)    <= sub_wire138(35);
	sub_wire2(119, 36)    <= sub_wire138(36);
	sub_wire2(119, 37)    <= sub_wire138(37);
	sub_wire2(119, 38)    <= sub_wire138(38);
	sub_wire2(119, 39)    <= sub_wire138(39);
	sub_wire2(118, 0)    <= sub_wire139(0);
	sub_wire2(118, 1)    <= sub_wire139(1);
	sub_wire2(118, 2)    <= sub_wire139(2);
	sub_wire2(118, 3)    <= sub_wire139(3);
	sub_wire2(118, 4)    <= sub_wire139(4);
	sub_wire2(118, 5)    <= sub_wire139(5);
	sub_wire2(118, 6)    <= sub_wire139(6);
	sub_wire2(118, 7)    <= sub_wire139(7);
	sub_wire2(118, 8)    <= sub_wire139(8);
	sub_wire2(118, 9)    <= sub_wire139(9);
	sub_wire2(118, 10)    <= sub_wire139(10);
	sub_wire2(118, 11)    <= sub_wire139(11);
	sub_wire2(118, 12)    <= sub_wire139(12);
	sub_wire2(118, 13)    <= sub_wire139(13);
	sub_wire2(118, 14)    <= sub_wire139(14);
	sub_wire2(118, 15)    <= sub_wire139(15);
	sub_wire2(118, 16)    <= sub_wire139(16);
	sub_wire2(118, 17)    <= sub_wire139(17);
	sub_wire2(118, 18)    <= sub_wire139(18);
	sub_wire2(118, 19)    <= sub_wire139(19);
	sub_wire2(118, 20)    <= sub_wire139(20);
	sub_wire2(118, 21)    <= sub_wire139(21);
	sub_wire2(118, 22)    <= sub_wire139(22);
	sub_wire2(118, 23)    <= sub_wire139(23);
	sub_wire2(118, 24)    <= sub_wire139(24);
	sub_wire2(118, 25)    <= sub_wire139(25);
	sub_wire2(118, 26)    <= sub_wire139(26);
	sub_wire2(118, 27)    <= sub_wire139(27);
	sub_wire2(118, 28)    <= sub_wire139(28);
	sub_wire2(118, 29)    <= sub_wire139(29);
	sub_wire2(118, 30)    <= sub_wire139(30);
	sub_wire2(118, 31)    <= sub_wire139(31);
	sub_wire2(118, 32)    <= sub_wire139(32);
	sub_wire2(118, 33)    <= sub_wire139(33);
	sub_wire2(118, 34)    <= sub_wire139(34);
	sub_wire2(118, 35)    <= sub_wire139(35);
	sub_wire2(118, 36)    <= sub_wire139(36);
	sub_wire2(118, 37)    <= sub_wire139(37);
	sub_wire2(118, 38)    <= sub_wire139(38);
	sub_wire2(118, 39)    <= sub_wire139(39);
	sub_wire2(117, 0)    <= sub_wire140(0);
	sub_wire2(117, 1)    <= sub_wire140(1);
	sub_wire2(117, 2)    <= sub_wire140(2);
	sub_wire2(117, 3)    <= sub_wire140(3);
	sub_wire2(117, 4)    <= sub_wire140(4);
	sub_wire2(117, 5)    <= sub_wire140(5);
	sub_wire2(117, 6)    <= sub_wire140(6);
	sub_wire2(117, 7)    <= sub_wire140(7);
	sub_wire2(117, 8)    <= sub_wire140(8);
	sub_wire2(117, 9)    <= sub_wire140(9);
	sub_wire2(117, 10)    <= sub_wire140(10);
	sub_wire2(117, 11)    <= sub_wire140(11);
	sub_wire2(117, 12)    <= sub_wire140(12);
	sub_wire2(117, 13)    <= sub_wire140(13);
	sub_wire2(117, 14)    <= sub_wire140(14);
	sub_wire2(117, 15)    <= sub_wire140(15);
	sub_wire2(117, 16)    <= sub_wire140(16);
	sub_wire2(117, 17)    <= sub_wire140(17);
	sub_wire2(117, 18)    <= sub_wire140(18);
	sub_wire2(117, 19)    <= sub_wire140(19);
	sub_wire2(117, 20)    <= sub_wire140(20);
	sub_wire2(117, 21)    <= sub_wire140(21);
	sub_wire2(117, 22)    <= sub_wire140(22);
	sub_wire2(117, 23)    <= sub_wire140(23);
	sub_wire2(117, 24)    <= sub_wire140(24);
	sub_wire2(117, 25)    <= sub_wire140(25);
	sub_wire2(117, 26)    <= sub_wire140(26);
	sub_wire2(117, 27)    <= sub_wire140(27);
	sub_wire2(117, 28)    <= sub_wire140(28);
	sub_wire2(117, 29)    <= sub_wire140(29);
	sub_wire2(117, 30)    <= sub_wire140(30);
	sub_wire2(117, 31)    <= sub_wire140(31);
	sub_wire2(117, 32)    <= sub_wire140(32);
	sub_wire2(117, 33)    <= sub_wire140(33);
	sub_wire2(117, 34)    <= sub_wire140(34);
	sub_wire2(117, 35)    <= sub_wire140(35);
	sub_wire2(117, 36)    <= sub_wire140(36);
	sub_wire2(117, 37)    <= sub_wire140(37);
	sub_wire2(117, 38)    <= sub_wire140(38);
	sub_wire2(117, 39)    <= sub_wire140(39);
	sub_wire2(116, 0)    <= sub_wire141(0);
	sub_wire2(116, 1)    <= sub_wire141(1);
	sub_wire2(116, 2)    <= sub_wire141(2);
	sub_wire2(116, 3)    <= sub_wire141(3);
	sub_wire2(116, 4)    <= sub_wire141(4);
	sub_wire2(116, 5)    <= sub_wire141(5);
	sub_wire2(116, 6)    <= sub_wire141(6);
	sub_wire2(116, 7)    <= sub_wire141(7);
	sub_wire2(116, 8)    <= sub_wire141(8);
	sub_wire2(116, 9)    <= sub_wire141(9);
	sub_wire2(116, 10)    <= sub_wire141(10);
	sub_wire2(116, 11)    <= sub_wire141(11);
	sub_wire2(116, 12)    <= sub_wire141(12);
	sub_wire2(116, 13)    <= sub_wire141(13);
	sub_wire2(116, 14)    <= sub_wire141(14);
	sub_wire2(116, 15)    <= sub_wire141(15);
	sub_wire2(116, 16)    <= sub_wire141(16);
	sub_wire2(116, 17)    <= sub_wire141(17);
	sub_wire2(116, 18)    <= sub_wire141(18);
	sub_wire2(116, 19)    <= sub_wire141(19);
	sub_wire2(116, 20)    <= sub_wire141(20);
	sub_wire2(116, 21)    <= sub_wire141(21);
	sub_wire2(116, 22)    <= sub_wire141(22);
	sub_wire2(116, 23)    <= sub_wire141(23);
	sub_wire2(116, 24)    <= sub_wire141(24);
	sub_wire2(116, 25)    <= sub_wire141(25);
	sub_wire2(116, 26)    <= sub_wire141(26);
	sub_wire2(116, 27)    <= sub_wire141(27);
	sub_wire2(116, 28)    <= sub_wire141(28);
	sub_wire2(116, 29)    <= sub_wire141(29);
	sub_wire2(116, 30)    <= sub_wire141(30);
	sub_wire2(116, 31)    <= sub_wire141(31);
	sub_wire2(116, 32)    <= sub_wire141(32);
	sub_wire2(116, 33)    <= sub_wire141(33);
	sub_wire2(116, 34)    <= sub_wire141(34);
	sub_wire2(116, 35)    <= sub_wire141(35);
	sub_wire2(116, 36)    <= sub_wire141(36);
	sub_wire2(116, 37)    <= sub_wire141(37);
	sub_wire2(116, 38)    <= sub_wire141(38);
	sub_wire2(116, 39)    <= sub_wire141(39);
	sub_wire2(115, 0)    <= sub_wire142(0);
	sub_wire2(115, 1)    <= sub_wire142(1);
	sub_wire2(115, 2)    <= sub_wire142(2);
	sub_wire2(115, 3)    <= sub_wire142(3);
	sub_wire2(115, 4)    <= sub_wire142(4);
	sub_wire2(115, 5)    <= sub_wire142(5);
	sub_wire2(115, 6)    <= sub_wire142(6);
	sub_wire2(115, 7)    <= sub_wire142(7);
	sub_wire2(115, 8)    <= sub_wire142(8);
	sub_wire2(115, 9)    <= sub_wire142(9);
	sub_wire2(115, 10)    <= sub_wire142(10);
	sub_wire2(115, 11)    <= sub_wire142(11);
	sub_wire2(115, 12)    <= sub_wire142(12);
	sub_wire2(115, 13)    <= sub_wire142(13);
	sub_wire2(115, 14)    <= sub_wire142(14);
	sub_wire2(115, 15)    <= sub_wire142(15);
	sub_wire2(115, 16)    <= sub_wire142(16);
	sub_wire2(115, 17)    <= sub_wire142(17);
	sub_wire2(115, 18)    <= sub_wire142(18);
	sub_wire2(115, 19)    <= sub_wire142(19);
	sub_wire2(115, 20)    <= sub_wire142(20);
	sub_wire2(115, 21)    <= sub_wire142(21);
	sub_wire2(115, 22)    <= sub_wire142(22);
	sub_wire2(115, 23)    <= sub_wire142(23);
	sub_wire2(115, 24)    <= sub_wire142(24);
	sub_wire2(115, 25)    <= sub_wire142(25);
	sub_wire2(115, 26)    <= sub_wire142(26);
	sub_wire2(115, 27)    <= sub_wire142(27);
	sub_wire2(115, 28)    <= sub_wire142(28);
	sub_wire2(115, 29)    <= sub_wire142(29);
	sub_wire2(115, 30)    <= sub_wire142(30);
	sub_wire2(115, 31)    <= sub_wire142(31);
	sub_wire2(115, 32)    <= sub_wire142(32);
	sub_wire2(115, 33)    <= sub_wire142(33);
	sub_wire2(115, 34)    <= sub_wire142(34);
	sub_wire2(115, 35)    <= sub_wire142(35);
	sub_wire2(115, 36)    <= sub_wire142(36);
	sub_wire2(115, 37)    <= sub_wire142(37);
	sub_wire2(115, 38)    <= sub_wire142(38);
	sub_wire2(115, 39)    <= sub_wire142(39);
	sub_wire2(114, 0)    <= sub_wire143(0);
	sub_wire2(114, 1)    <= sub_wire143(1);
	sub_wire2(114, 2)    <= sub_wire143(2);
	sub_wire2(114, 3)    <= sub_wire143(3);
	sub_wire2(114, 4)    <= sub_wire143(4);
	sub_wire2(114, 5)    <= sub_wire143(5);
	sub_wire2(114, 6)    <= sub_wire143(6);
	sub_wire2(114, 7)    <= sub_wire143(7);
	sub_wire2(114, 8)    <= sub_wire143(8);
	sub_wire2(114, 9)    <= sub_wire143(9);
	sub_wire2(114, 10)    <= sub_wire143(10);
	sub_wire2(114, 11)    <= sub_wire143(11);
	sub_wire2(114, 12)    <= sub_wire143(12);
	sub_wire2(114, 13)    <= sub_wire143(13);
	sub_wire2(114, 14)    <= sub_wire143(14);
	sub_wire2(114, 15)    <= sub_wire143(15);
	sub_wire2(114, 16)    <= sub_wire143(16);
	sub_wire2(114, 17)    <= sub_wire143(17);
	sub_wire2(114, 18)    <= sub_wire143(18);
	sub_wire2(114, 19)    <= sub_wire143(19);
	sub_wire2(114, 20)    <= sub_wire143(20);
	sub_wire2(114, 21)    <= sub_wire143(21);
	sub_wire2(114, 22)    <= sub_wire143(22);
	sub_wire2(114, 23)    <= sub_wire143(23);
	sub_wire2(114, 24)    <= sub_wire143(24);
	sub_wire2(114, 25)    <= sub_wire143(25);
	sub_wire2(114, 26)    <= sub_wire143(26);
	sub_wire2(114, 27)    <= sub_wire143(27);
	sub_wire2(114, 28)    <= sub_wire143(28);
	sub_wire2(114, 29)    <= sub_wire143(29);
	sub_wire2(114, 30)    <= sub_wire143(30);
	sub_wire2(114, 31)    <= sub_wire143(31);
	sub_wire2(114, 32)    <= sub_wire143(32);
	sub_wire2(114, 33)    <= sub_wire143(33);
	sub_wire2(114, 34)    <= sub_wire143(34);
	sub_wire2(114, 35)    <= sub_wire143(35);
	sub_wire2(114, 36)    <= sub_wire143(36);
	sub_wire2(114, 37)    <= sub_wire143(37);
	sub_wire2(114, 38)    <= sub_wire143(38);
	sub_wire2(114, 39)    <= sub_wire143(39);
	sub_wire2(113, 0)    <= sub_wire144(0);
	sub_wire2(113, 1)    <= sub_wire144(1);
	sub_wire2(113, 2)    <= sub_wire144(2);
	sub_wire2(113, 3)    <= sub_wire144(3);
	sub_wire2(113, 4)    <= sub_wire144(4);
	sub_wire2(113, 5)    <= sub_wire144(5);
	sub_wire2(113, 6)    <= sub_wire144(6);
	sub_wire2(113, 7)    <= sub_wire144(7);
	sub_wire2(113, 8)    <= sub_wire144(8);
	sub_wire2(113, 9)    <= sub_wire144(9);
	sub_wire2(113, 10)    <= sub_wire144(10);
	sub_wire2(113, 11)    <= sub_wire144(11);
	sub_wire2(113, 12)    <= sub_wire144(12);
	sub_wire2(113, 13)    <= sub_wire144(13);
	sub_wire2(113, 14)    <= sub_wire144(14);
	sub_wire2(113, 15)    <= sub_wire144(15);
	sub_wire2(113, 16)    <= sub_wire144(16);
	sub_wire2(113, 17)    <= sub_wire144(17);
	sub_wire2(113, 18)    <= sub_wire144(18);
	sub_wire2(113, 19)    <= sub_wire144(19);
	sub_wire2(113, 20)    <= sub_wire144(20);
	sub_wire2(113, 21)    <= sub_wire144(21);
	sub_wire2(113, 22)    <= sub_wire144(22);
	sub_wire2(113, 23)    <= sub_wire144(23);
	sub_wire2(113, 24)    <= sub_wire144(24);
	sub_wire2(113, 25)    <= sub_wire144(25);
	sub_wire2(113, 26)    <= sub_wire144(26);
	sub_wire2(113, 27)    <= sub_wire144(27);
	sub_wire2(113, 28)    <= sub_wire144(28);
	sub_wire2(113, 29)    <= sub_wire144(29);
	sub_wire2(113, 30)    <= sub_wire144(30);
	sub_wire2(113, 31)    <= sub_wire144(31);
	sub_wire2(113, 32)    <= sub_wire144(32);
	sub_wire2(113, 33)    <= sub_wire144(33);
	sub_wire2(113, 34)    <= sub_wire144(34);
	sub_wire2(113, 35)    <= sub_wire144(35);
	sub_wire2(113, 36)    <= sub_wire144(36);
	sub_wire2(113, 37)    <= sub_wire144(37);
	sub_wire2(113, 38)    <= sub_wire144(38);
	sub_wire2(113, 39)    <= sub_wire144(39);
	sub_wire2(112, 0)    <= sub_wire145(0);
	sub_wire2(112, 1)    <= sub_wire145(1);
	sub_wire2(112, 2)    <= sub_wire145(2);
	sub_wire2(112, 3)    <= sub_wire145(3);
	sub_wire2(112, 4)    <= sub_wire145(4);
	sub_wire2(112, 5)    <= sub_wire145(5);
	sub_wire2(112, 6)    <= sub_wire145(6);
	sub_wire2(112, 7)    <= sub_wire145(7);
	sub_wire2(112, 8)    <= sub_wire145(8);
	sub_wire2(112, 9)    <= sub_wire145(9);
	sub_wire2(112, 10)    <= sub_wire145(10);
	sub_wire2(112, 11)    <= sub_wire145(11);
	sub_wire2(112, 12)    <= sub_wire145(12);
	sub_wire2(112, 13)    <= sub_wire145(13);
	sub_wire2(112, 14)    <= sub_wire145(14);
	sub_wire2(112, 15)    <= sub_wire145(15);
	sub_wire2(112, 16)    <= sub_wire145(16);
	sub_wire2(112, 17)    <= sub_wire145(17);
	sub_wire2(112, 18)    <= sub_wire145(18);
	sub_wire2(112, 19)    <= sub_wire145(19);
	sub_wire2(112, 20)    <= sub_wire145(20);
	sub_wire2(112, 21)    <= sub_wire145(21);
	sub_wire2(112, 22)    <= sub_wire145(22);
	sub_wire2(112, 23)    <= sub_wire145(23);
	sub_wire2(112, 24)    <= sub_wire145(24);
	sub_wire2(112, 25)    <= sub_wire145(25);
	sub_wire2(112, 26)    <= sub_wire145(26);
	sub_wire2(112, 27)    <= sub_wire145(27);
	sub_wire2(112, 28)    <= sub_wire145(28);
	sub_wire2(112, 29)    <= sub_wire145(29);
	sub_wire2(112, 30)    <= sub_wire145(30);
	sub_wire2(112, 31)    <= sub_wire145(31);
	sub_wire2(112, 32)    <= sub_wire145(32);
	sub_wire2(112, 33)    <= sub_wire145(33);
	sub_wire2(112, 34)    <= sub_wire145(34);
	sub_wire2(112, 35)    <= sub_wire145(35);
	sub_wire2(112, 36)    <= sub_wire145(36);
	sub_wire2(112, 37)    <= sub_wire145(37);
	sub_wire2(112, 38)    <= sub_wire145(38);
	sub_wire2(112, 39)    <= sub_wire145(39);
	sub_wire2(111, 0)    <= sub_wire146(0);
	sub_wire2(111, 1)    <= sub_wire146(1);
	sub_wire2(111, 2)    <= sub_wire146(2);
	sub_wire2(111, 3)    <= sub_wire146(3);
	sub_wire2(111, 4)    <= sub_wire146(4);
	sub_wire2(111, 5)    <= sub_wire146(5);
	sub_wire2(111, 6)    <= sub_wire146(6);
	sub_wire2(111, 7)    <= sub_wire146(7);
	sub_wire2(111, 8)    <= sub_wire146(8);
	sub_wire2(111, 9)    <= sub_wire146(9);
	sub_wire2(111, 10)    <= sub_wire146(10);
	sub_wire2(111, 11)    <= sub_wire146(11);
	sub_wire2(111, 12)    <= sub_wire146(12);
	sub_wire2(111, 13)    <= sub_wire146(13);
	sub_wire2(111, 14)    <= sub_wire146(14);
	sub_wire2(111, 15)    <= sub_wire146(15);
	sub_wire2(111, 16)    <= sub_wire146(16);
	sub_wire2(111, 17)    <= sub_wire146(17);
	sub_wire2(111, 18)    <= sub_wire146(18);
	sub_wire2(111, 19)    <= sub_wire146(19);
	sub_wire2(111, 20)    <= sub_wire146(20);
	sub_wire2(111, 21)    <= sub_wire146(21);
	sub_wire2(111, 22)    <= sub_wire146(22);
	sub_wire2(111, 23)    <= sub_wire146(23);
	sub_wire2(111, 24)    <= sub_wire146(24);
	sub_wire2(111, 25)    <= sub_wire146(25);
	sub_wire2(111, 26)    <= sub_wire146(26);
	sub_wire2(111, 27)    <= sub_wire146(27);
	sub_wire2(111, 28)    <= sub_wire146(28);
	sub_wire2(111, 29)    <= sub_wire146(29);
	sub_wire2(111, 30)    <= sub_wire146(30);
	sub_wire2(111, 31)    <= sub_wire146(31);
	sub_wire2(111, 32)    <= sub_wire146(32);
	sub_wire2(111, 33)    <= sub_wire146(33);
	sub_wire2(111, 34)    <= sub_wire146(34);
	sub_wire2(111, 35)    <= sub_wire146(35);
	sub_wire2(111, 36)    <= sub_wire146(36);
	sub_wire2(111, 37)    <= sub_wire146(37);
	sub_wire2(111, 38)    <= sub_wire146(38);
	sub_wire2(111, 39)    <= sub_wire146(39);
	sub_wire2(110, 0)    <= sub_wire147(0);
	sub_wire2(110, 1)    <= sub_wire147(1);
	sub_wire2(110, 2)    <= sub_wire147(2);
	sub_wire2(110, 3)    <= sub_wire147(3);
	sub_wire2(110, 4)    <= sub_wire147(4);
	sub_wire2(110, 5)    <= sub_wire147(5);
	sub_wire2(110, 6)    <= sub_wire147(6);
	sub_wire2(110, 7)    <= sub_wire147(7);
	sub_wire2(110, 8)    <= sub_wire147(8);
	sub_wire2(110, 9)    <= sub_wire147(9);
	sub_wire2(110, 10)    <= sub_wire147(10);
	sub_wire2(110, 11)    <= sub_wire147(11);
	sub_wire2(110, 12)    <= sub_wire147(12);
	sub_wire2(110, 13)    <= sub_wire147(13);
	sub_wire2(110, 14)    <= sub_wire147(14);
	sub_wire2(110, 15)    <= sub_wire147(15);
	sub_wire2(110, 16)    <= sub_wire147(16);
	sub_wire2(110, 17)    <= sub_wire147(17);
	sub_wire2(110, 18)    <= sub_wire147(18);
	sub_wire2(110, 19)    <= sub_wire147(19);
	sub_wire2(110, 20)    <= sub_wire147(20);
	sub_wire2(110, 21)    <= sub_wire147(21);
	sub_wire2(110, 22)    <= sub_wire147(22);
	sub_wire2(110, 23)    <= sub_wire147(23);
	sub_wire2(110, 24)    <= sub_wire147(24);
	sub_wire2(110, 25)    <= sub_wire147(25);
	sub_wire2(110, 26)    <= sub_wire147(26);
	sub_wire2(110, 27)    <= sub_wire147(27);
	sub_wire2(110, 28)    <= sub_wire147(28);
	sub_wire2(110, 29)    <= sub_wire147(29);
	sub_wire2(110, 30)    <= sub_wire147(30);
	sub_wire2(110, 31)    <= sub_wire147(31);
	sub_wire2(110, 32)    <= sub_wire147(32);
	sub_wire2(110, 33)    <= sub_wire147(33);
	sub_wire2(110, 34)    <= sub_wire147(34);
	sub_wire2(110, 35)    <= sub_wire147(35);
	sub_wire2(110, 36)    <= sub_wire147(36);
	sub_wire2(110, 37)    <= sub_wire147(37);
	sub_wire2(110, 38)    <= sub_wire147(38);
	sub_wire2(110, 39)    <= sub_wire147(39);
	sub_wire2(109, 0)    <= sub_wire148(0);
	sub_wire2(109, 1)    <= sub_wire148(1);
	sub_wire2(109, 2)    <= sub_wire148(2);
	sub_wire2(109, 3)    <= sub_wire148(3);
	sub_wire2(109, 4)    <= sub_wire148(4);
	sub_wire2(109, 5)    <= sub_wire148(5);
	sub_wire2(109, 6)    <= sub_wire148(6);
	sub_wire2(109, 7)    <= sub_wire148(7);
	sub_wire2(109, 8)    <= sub_wire148(8);
	sub_wire2(109, 9)    <= sub_wire148(9);
	sub_wire2(109, 10)    <= sub_wire148(10);
	sub_wire2(109, 11)    <= sub_wire148(11);
	sub_wire2(109, 12)    <= sub_wire148(12);
	sub_wire2(109, 13)    <= sub_wire148(13);
	sub_wire2(109, 14)    <= sub_wire148(14);
	sub_wire2(109, 15)    <= sub_wire148(15);
	sub_wire2(109, 16)    <= sub_wire148(16);
	sub_wire2(109, 17)    <= sub_wire148(17);
	sub_wire2(109, 18)    <= sub_wire148(18);
	sub_wire2(109, 19)    <= sub_wire148(19);
	sub_wire2(109, 20)    <= sub_wire148(20);
	sub_wire2(109, 21)    <= sub_wire148(21);
	sub_wire2(109, 22)    <= sub_wire148(22);
	sub_wire2(109, 23)    <= sub_wire148(23);
	sub_wire2(109, 24)    <= sub_wire148(24);
	sub_wire2(109, 25)    <= sub_wire148(25);
	sub_wire2(109, 26)    <= sub_wire148(26);
	sub_wire2(109, 27)    <= sub_wire148(27);
	sub_wire2(109, 28)    <= sub_wire148(28);
	sub_wire2(109, 29)    <= sub_wire148(29);
	sub_wire2(109, 30)    <= sub_wire148(30);
	sub_wire2(109, 31)    <= sub_wire148(31);
	sub_wire2(109, 32)    <= sub_wire148(32);
	sub_wire2(109, 33)    <= sub_wire148(33);
	sub_wire2(109, 34)    <= sub_wire148(34);
	sub_wire2(109, 35)    <= sub_wire148(35);
	sub_wire2(109, 36)    <= sub_wire148(36);
	sub_wire2(109, 37)    <= sub_wire148(37);
	sub_wire2(109, 38)    <= sub_wire148(38);
	sub_wire2(109, 39)    <= sub_wire148(39);
	sub_wire2(108, 0)    <= sub_wire149(0);
	sub_wire2(108, 1)    <= sub_wire149(1);
	sub_wire2(108, 2)    <= sub_wire149(2);
	sub_wire2(108, 3)    <= sub_wire149(3);
	sub_wire2(108, 4)    <= sub_wire149(4);
	sub_wire2(108, 5)    <= sub_wire149(5);
	sub_wire2(108, 6)    <= sub_wire149(6);
	sub_wire2(108, 7)    <= sub_wire149(7);
	sub_wire2(108, 8)    <= sub_wire149(8);
	sub_wire2(108, 9)    <= sub_wire149(9);
	sub_wire2(108, 10)    <= sub_wire149(10);
	sub_wire2(108, 11)    <= sub_wire149(11);
	sub_wire2(108, 12)    <= sub_wire149(12);
	sub_wire2(108, 13)    <= sub_wire149(13);
	sub_wire2(108, 14)    <= sub_wire149(14);
	sub_wire2(108, 15)    <= sub_wire149(15);
	sub_wire2(108, 16)    <= sub_wire149(16);
	sub_wire2(108, 17)    <= sub_wire149(17);
	sub_wire2(108, 18)    <= sub_wire149(18);
	sub_wire2(108, 19)    <= sub_wire149(19);
	sub_wire2(108, 20)    <= sub_wire149(20);
	sub_wire2(108, 21)    <= sub_wire149(21);
	sub_wire2(108, 22)    <= sub_wire149(22);
	sub_wire2(108, 23)    <= sub_wire149(23);
	sub_wire2(108, 24)    <= sub_wire149(24);
	sub_wire2(108, 25)    <= sub_wire149(25);
	sub_wire2(108, 26)    <= sub_wire149(26);
	sub_wire2(108, 27)    <= sub_wire149(27);
	sub_wire2(108, 28)    <= sub_wire149(28);
	sub_wire2(108, 29)    <= sub_wire149(29);
	sub_wire2(108, 30)    <= sub_wire149(30);
	sub_wire2(108, 31)    <= sub_wire149(31);
	sub_wire2(108, 32)    <= sub_wire149(32);
	sub_wire2(108, 33)    <= sub_wire149(33);
	sub_wire2(108, 34)    <= sub_wire149(34);
	sub_wire2(108, 35)    <= sub_wire149(35);
	sub_wire2(108, 36)    <= sub_wire149(36);
	sub_wire2(108, 37)    <= sub_wire149(37);
	sub_wire2(108, 38)    <= sub_wire149(38);
	sub_wire2(108, 39)    <= sub_wire149(39);
	sub_wire2(107, 0)    <= sub_wire150(0);
	sub_wire2(107, 1)    <= sub_wire150(1);
	sub_wire2(107, 2)    <= sub_wire150(2);
	sub_wire2(107, 3)    <= sub_wire150(3);
	sub_wire2(107, 4)    <= sub_wire150(4);
	sub_wire2(107, 5)    <= sub_wire150(5);
	sub_wire2(107, 6)    <= sub_wire150(6);
	sub_wire2(107, 7)    <= sub_wire150(7);
	sub_wire2(107, 8)    <= sub_wire150(8);
	sub_wire2(107, 9)    <= sub_wire150(9);
	sub_wire2(107, 10)    <= sub_wire150(10);
	sub_wire2(107, 11)    <= sub_wire150(11);
	sub_wire2(107, 12)    <= sub_wire150(12);
	sub_wire2(107, 13)    <= sub_wire150(13);
	sub_wire2(107, 14)    <= sub_wire150(14);
	sub_wire2(107, 15)    <= sub_wire150(15);
	sub_wire2(107, 16)    <= sub_wire150(16);
	sub_wire2(107, 17)    <= sub_wire150(17);
	sub_wire2(107, 18)    <= sub_wire150(18);
	sub_wire2(107, 19)    <= sub_wire150(19);
	sub_wire2(107, 20)    <= sub_wire150(20);
	sub_wire2(107, 21)    <= sub_wire150(21);
	sub_wire2(107, 22)    <= sub_wire150(22);
	sub_wire2(107, 23)    <= sub_wire150(23);
	sub_wire2(107, 24)    <= sub_wire150(24);
	sub_wire2(107, 25)    <= sub_wire150(25);
	sub_wire2(107, 26)    <= sub_wire150(26);
	sub_wire2(107, 27)    <= sub_wire150(27);
	sub_wire2(107, 28)    <= sub_wire150(28);
	sub_wire2(107, 29)    <= sub_wire150(29);
	sub_wire2(107, 30)    <= sub_wire150(30);
	sub_wire2(107, 31)    <= sub_wire150(31);
	sub_wire2(107, 32)    <= sub_wire150(32);
	sub_wire2(107, 33)    <= sub_wire150(33);
	sub_wire2(107, 34)    <= sub_wire150(34);
	sub_wire2(107, 35)    <= sub_wire150(35);
	sub_wire2(107, 36)    <= sub_wire150(36);
	sub_wire2(107, 37)    <= sub_wire150(37);
	sub_wire2(107, 38)    <= sub_wire150(38);
	sub_wire2(107, 39)    <= sub_wire150(39);
	sub_wire2(106, 0)    <= sub_wire151(0);
	sub_wire2(106, 1)    <= sub_wire151(1);
	sub_wire2(106, 2)    <= sub_wire151(2);
	sub_wire2(106, 3)    <= sub_wire151(3);
	sub_wire2(106, 4)    <= sub_wire151(4);
	sub_wire2(106, 5)    <= sub_wire151(5);
	sub_wire2(106, 6)    <= sub_wire151(6);
	sub_wire2(106, 7)    <= sub_wire151(7);
	sub_wire2(106, 8)    <= sub_wire151(8);
	sub_wire2(106, 9)    <= sub_wire151(9);
	sub_wire2(106, 10)    <= sub_wire151(10);
	sub_wire2(106, 11)    <= sub_wire151(11);
	sub_wire2(106, 12)    <= sub_wire151(12);
	sub_wire2(106, 13)    <= sub_wire151(13);
	sub_wire2(106, 14)    <= sub_wire151(14);
	sub_wire2(106, 15)    <= sub_wire151(15);
	sub_wire2(106, 16)    <= sub_wire151(16);
	sub_wire2(106, 17)    <= sub_wire151(17);
	sub_wire2(106, 18)    <= sub_wire151(18);
	sub_wire2(106, 19)    <= sub_wire151(19);
	sub_wire2(106, 20)    <= sub_wire151(20);
	sub_wire2(106, 21)    <= sub_wire151(21);
	sub_wire2(106, 22)    <= sub_wire151(22);
	sub_wire2(106, 23)    <= sub_wire151(23);
	sub_wire2(106, 24)    <= sub_wire151(24);
	sub_wire2(106, 25)    <= sub_wire151(25);
	sub_wire2(106, 26)    <= sub_wire151(26);
	sub_wire2(106, 27)    <= sub_wire151(27);
	sub_wire2(106, 28)    <= sub_wire151(28);
	sub_wire2(106, 29)    <= sub_wire151(29);
	sub_wire2(106, 30)    <= sub_wire151(30);
	sub_wire2(106, 31)    <= sub_wire151(31);
	sub_wire2(106, 32)    <= sub_wire151(32);
	sub_wire2(106, 33)    <= sub_wire151(33);
	sub_wire2(106, 34)    <= sub_wire151(34);
	sub_wire2(106, 35)    <= sub_wire151(35);
	sub_wire2(106, 36)    <= sub_wire151(36);
	sub_wire2(106, 37)    <= sub_wire151(37);
	sub_wire2(106, 38)    <= sub_wire151(38);
	sub_wire2(106, 39)    <= sub_wire151(39);
	sub_wire2(105, 0)    <= sub_wire152(0);
	sub_wire2(105, 1)    <= sub_wire152(1);
	sub_wire2(105, 2)    <= sub_wire152(2);
	sub_wire2(105, 3)    <= sub_wire152(3);
	sub_wire2(105, 4)    <= sub_wire152(4);
	sub_wire2(105, 5)    <= sub_wire152(5);
	sub_wire2(105, 6)    <= sub_wire152(6);
	sub_wire2(105, 7)    <= sub_wire152(7);
	sub_wire2(105, 8)    <= sub_wire152(8);
	sub_wire2(105, 9)    <= sub_wire152(9);
	sub_wire2(105, 10)    <= sub_wire152(10);
	sub_wire2(105, 11)    <= sub_wire152(11);
	sub_wire2(105, 12)    <= sub_wire152(12);
	sub_wire2(105, 13)    <= sub_wire152(13);
	sub_wire2(105, 14)    <= sub_wire152(14);
	sub_wire2(105, 15)    <= sub_wire152(15);
	sub_wire2(105, 16)    <= sub_wire152(16);
	sub_wire2(105, 17)    <= sub_wire152(17);
	sub_wire2(105, 18)    <= sub_wire152(18);
	sub_wire2(105, 19)    <= sub_wire152(19);
	sub_wire2(105, 20)    <= sub_wire152(20);
	sub_wire2(105, 21)    <= sub_wire152(21);
	sub_wire2(105, 22)    <= sub_wire152(22);
	sub_wire2(105, 23)    <= sub_wire152(23);
	sub_wire2(105, 24)    <= sub_wire152(24);
	sub_wire2(105, 25)    <= sub_wire152(25);
	sub_wire2(105, 26)    <= sub_wire152(26);
	sub_wire2(105, 27)    <= sub_wire152(27);
	sub_wire2(105, 28)    <= sub_wire152(28);
	sub_wire2(105, 29)    <= sub_wire152(29);
	sub_wire2(105, 30)    <= sub_wire152(30);
	sub_wire2(105, 31)    <= sub_wire152(31);
	sub_wire2(105, 32)    <= sub_wire152(32);
	sub_wire2(105, 33)    <= sub_wire152(33);
	sub_wire2(105, 34)    <= sub_wire152(34);
	sub_wire2(105, 35)    <= sub_wire152(35);
	sub_wire2(105, 36)    <= sub_wire152(36);
	sub_wire2(105, 37)    <= sub_wire152(37);
	sub_wire2(105, 38)    <= sub_wire152(38);
	sub_wire2(105, 39)    <= sub_wire152(39);
	sub_wire2(104, 0)    <= sub_wire153(0);
	sub_wire2(104, 1)    <= sub_wire153(1);
	sub_wire2(104, 2)    <= sub_wire153(2);
	sub_wire2(104, 3)    <= sub_wire153(3);
	sub_wire2(104, 4)    <= sub_wire153(4);
	sub_wire2(104, 5)    <= sub_wire153(5);
	sub_wire2(104, 6)    <= sub_wire153(6);
	sub_wire2(104, 7)    <= sub_wire153(7);
	sub_wire2(104, 8)    <= sub_wire153(8);
	sub_wire2(104, 9)    <= sub_wire153(9);
	sub_wire2(104, 10)    <= sub_wire153(10);
	sub_wire2(104, 11)    <= sub_wire153(11);
	sub_wire2(104, 12)    <= sub_wire153(12);
	sub_wire2(104, 13)    <= sub_wire153(13);
	sub_wire2(104, 14)    <= sub_wire153(14);
	sub_wire2(104, 15)    <= sub_wire153(15);
	sub_wire2(104, 16)    <= sub_wire153(16);
	sub_wire2(104, 17)    <= sub_wire153(17);
	sub_wire2(104, 18)    <= sub_wire153(18);
	sub_wire2(104, 19)    <= sub_wire153(19);
	sub_wire2(104, 20)    <= sub_wire153(20);
	sub_wire2(104, 21)    <= sub_wire153(21);
	sub_wire2(104, 22)    <= sub_wire153(22);
	sub_wire2(104, 23)    <= sub_wire153(23);
	sub_wire2(104, 24)    <= sub_wire153(24);
	sub_wire2(104, 25)    <= sub_wire153(25);
	sub_wire2(104, 26)    <= sub_wire153(26);
	sub_wire2(104, 27)    <= sub_wire153(27);
	sub_wire2(104, 28)    <= sub_wire153(28);
	sub_wire2(104, 29)    <= sub_wire153(29);
	sub_wire2(104, 30)    <= sub_wire153(30);
	sub_wire2(104, 31)    <= sub_wire153(31);
	sub_wire2(104, 32)    <= sub_wire153(32);
	sub_wire2(104, 33)    <= sub_wire153(33);
	sub_wire2(104, 34)    <= sub_wire153(34);
	sub_wire2(104, 35)    <= sub_wire153(35);
	sub_wire2(104, 36)    <= sub_wire153(36);
	sub_wire2(104, 37)    <= sub_wire153(37);
	sub_wire2(104, 38)    <= sub_wire153(38);
	sub_wire2(104, 39)    <= sub_wire153(39);
	sub_wire2(103, 0)    <= sub_wire154(0);
	sub_wire2(103, 1)    <= sub_wire154(1);
	sub_wire2(103, 2)    <= sub_wire154(2);
	sub_wire2(103, 3)    <= sub_wire154(3);
	sub_wire2(103, 4)    <= sub_wire154(4);
	sub_wire2(103, 5)    <= sub_wire154(5);
	sub_wire2(103, 6)    <= sub_wire154(6);
	sub_wire2(103, 7)    <= sub_wire154(7);
	sub_wire2(103, 8)    <= sub_wire154(8);
	sub_wire2(103, 9)    <= sub_wire154(9);
	sub_wire2(103, 10)    <= sub_wire154(10);
	sub_wire2(103, 11)    <= sub_wire154(11);
	sub_wire2(103, 12)    <= sub_wire154(12);
	sub_wire2(103, 13)    <= sub_wire154(13);
	sub_wire2(103, 14)    <= sub_wire154(14);
	sub_wire2(103, 15)    <= sub_wire154(15);
	sub_wire2(103, 16)    <= sub_wire154(16);
	sub_wire2(103, 17)    <= sub_wire154(17);
	sub_wire2(103, 18)    <= sub_wire154(18);
	sub_wire2(103, 19)    <= sub_wire154(19);
	sub_wire2(103, 20)    <= sub_wire154(20);
	sub_wire2(103, 21)    <= sub_wire154(21);
	sub_wire2(103, 22)    <= sub_wire154(22);
	sub_wire2(103, 23)    <= sub_wire154(23);
	sub_wire2(103, 24)    <= sub_wire154(24);
	sub_wire2(103, 25)    <= sub_wire154(25);
	sub_wire2(103, 26)    <= sub_wire154(26);
	sub_wire2(103, 27)    <= sub_wire154(27);
	sub_wire2(103, 28)    <= sub_wire154(28);
	sub_wire2(103, 29)    <= sub_wire154(29);
	sub_wire2(103, 30)    <= sub_wire154(30);
	sub_wire2(103, 31)    <= sub_wire154(31);
	sub_wire2(103, 32)    <= sub_wire154(32);
	sub_wire2(103, 33)    <= sub_wire154(33);
	sub_wire2(103, 34)    <= sub_wire154(34);
	sub_wire2(103, 35)    <= sub_wire154(35);
	sub_wire2(103, 36)    <= sub_wire154(36);
	sub_wire2(103, 37)    <= sub_wire154(37);
	sub_wire2(103, 38)    <= sub_wire154(38);
	sub_wire2(103, 39)    <= sub_wire154(39);
	sub_wire2(102, 0)    <= sub_wire155(0);
	sub_wire2(102, 1)    <= sub_wire155(1);
	sub_wire2(102, 2)    <= sub_wire155(2);
	sub_wire2(102, 3)    <= sub_wire155(3);
	sub_wire2(102, 4)    <= sub_wire155(4);
	sub_wire2(102, 5)    <= sub_wire155(5);
	sub_wire2(102, 6)    <= sub_wire155(6);
	sub_wire2(102, 7)    <= sub_wire155(7);
	sub_wire2(102, 8)    <= sub_wire155(8);
	sub_wire2(102, 9)    <= sub_wire155(9);
	sub_wire2(102, 10)    <= sub_wire155(10);
	sub_wire2(102, 11)    <= sub_wire155(11);
	sub_wire2(102, 12)    <= sub_wire155(12);
	sub_wire2(102, 13)    <= sub_wire155(13);
	sub_wire2(102, 14)    <= sub_wire155(14);
	sub_wire2(102, 15)    <= sub_wire155(15);
	sub_wire2(102, 16)    <= sub_wire155(16);
	sub_wire2(102, 17)    <= sub_wire155(17);
	sub_wire2(102, 18)    <= sub_wire155(18);
	sub_wire2(102, 19)    <= sub_wire155(19);
	sub_wire2(102, 20)    <= sub_wire155(20);
	sub_wire2(102, 21)    <= sub_wire155(21);
	sub_wire2(102, 22)    <= sub_wire155(22);
	sub_wire2(102, 23)    <= sub_wire155(23);
	sub_wire2(102, 24)    <= sub_wire155(24);
	sub_wire2(102, 25)    <= sub_wire155(25);
	sub_wire2(102, 26)    <= sub_wire155(26);
	sub_wire2(102, 27)    <= sub_wire155(27);
	sub_wire2(102, 28)    <= sub_wire155(28);
	sub_wire2(102, 29)    <= sub_wire155(29);
	sub_wire2(102, 30)    <= sub_wire155(30);
	sub_wire2(102, 31)    <= sub_wire155(31);
	sub_wire2(102, 32)    <= sub_wire155(32);
	sub_wire2(102, 33)    <= sub_wire155(33);
	sub_wire2(102, 34)    <= sub_wire155(34);
	sub_wire2(102, 35)    <= sub_wire155(35);
	sub_wire2(102, 36)    <= sub_wire155(36);
	sub_wire2(102, 37)    <= sub_wire155(37);
	sub_wire2(102, 38)    <= sub_wire155(38);
	sub_wire2(102, 39)    <= sub_wire155(39);
	sub_wire2(101, 0)    <= sub_wire156(0);
	sub_wire2(101, 1)    <= sub_wire156(1);
	sub_wire2(101, 2)    <= sub_wire156(2);
	sub_wire2(101, 3)    <= sub_wire156(3);
	sub_wire2(101, 4)    <= sub_wire156(4);
	sub_wire2(101, 5)    <= sub_wire156(5);
	sub_wire2(101, 6)    <= sub_wire156(6);
	sub_wire2(101, 7)    <= sub_wire156(7);
	sub_wire2(101, 8)    <= sub_wire156(8);
	sub_wire2(101, 9)    <= sub_wire156(9);
	sub_wire2(101, 10)    <= sub_wire156(10);
	sub_wire2(101, 11)    <= sub_wire156(11);
	sub_wire2(101, 12)    <= sub_wire156(12);
	sub_wire2(101, 13)    <= sub_wire156(13);
	sub_wire2(101, 14)    <= sub_wire156(14);
	sub_wire2(101, 15)    <= sub_wire156(15);
	sub_wire2(101, 16)    <= sub_wire156(16);
	sub_wire2(101, 17)    <= sub_wire156(17);
	sub_wire2(101, 18)    <= sub_wire156(18);
	sub_wire2(101, 19)    <= sub_wire156(19);
	sub_wire2(101, 20)    <= sub_wire156(20);
	sub_wire2(101, 21)    <= sub_wire156(21);
	sub_wire2(101, 22)    <= sub_wire156(22);
	sub_wire2(101, 23)    <= sub_wire156(23);
	sub_wire2(101, 24)    <= sub_wire156(24);
	sub_wire2(101, 25)    <= sub_wire156(25);
	sub_wire2(101, 26)    <= sub_wire156(26);
	sub_wire2(101, 27)    <= sub_wire156(27);
	sub_wire2(101, 28)    <= sub_wire156(28);
	sub_wire2(101, 29)    <= sub_wire156(29);
	sub_wire2(101, 30)    <= sub_wire156(30);
	sub_wire2(101, 31)    <= sub_wire156(31);
	sub_wire2(101, 32)    <= sub_wire156(32);
	sub_wire2(101, 33)    <= sub_wire156(33);
	sub_wire2(101, 34)    <= sub_wire156(34);
	sub_wire2(101, 35)    <= sub_wire156(35);
	sub_wire2(101, 36)    <= sub_wire156(36);
	sub_wire2(101, 37)    <= sub_wire156(37);
	sub_wire2(101, 38)    <= sub_wire156(38);
	sub_wire2(101, 39)    <= sub_wire156(39);
	sub_wire2(100, 0)    <= sub_wire157(0);
	sub_wire2(100, 1)    <= sub_wire157(1);
	sub_wire2(100, 2)    <= sub_wire157(2);
	sub_wire2(100, 3)    <= sub_wire157(3);
	sub_wire2(100, 4)    <= sub_wire157(4);
	sub_wire2(100, 5)    <= sub_wire157(5);
	sub_wire2(100, 6)    <= sub_wire157(6);
	sub_wire2(100, 7)    <= sub_wire157(7);
	sub_wire2(100, 8)    <= sub_wire157(8);
	sub_wire2(100, 9)    <= sub_wire157(9);
	sub_wire2(100, 10)    <= sub_wire157(10);
	sub_wire2(100, 11)    <= sub_wire157(11);
	sub_wire2(100, 12)    <= sub_wire157(12);
	sub_wire2(100, 13)    <= sub_wire157(13);
	sub_wire2(100, 14)    <= sub_wire157(14);
	sub_wire2(100, 15)    <= sub_wire157(15);
	sub_wire2(100, 16)    <= sub_wire157(16);
	sub_wire2(100, 17)    <= sub_wire157(17);
	sub_wire2(100, 18)    <= sub_wire157(18);
	sub_wire2(100, 19)    <= sub_wire157(19);
	sub_wire2(100, 20)    <= sub_wire157(20);
	sub_wire2(100, 21)    <= sub_wire157(21);
	sub_wire2(100, 22)    <= sub_wire157(22);
	sub_wire2(100, 23)    <= sub_wire157(23);
	sub_wire2(100, 24)    <= sub_wire157(24);
	sub_wire2(100, 25)    <= sub_wire157(25);
	sub_wire2(100, 26)    <= sub_wire157(26);
	sub_wire2(100, 27)    <= sub_wire157(27);
	sub_wire2(100, 28)    <= sub_wire157(28);
	sub_wire2(100, 29)    <= sub_wire157(29);
	sub_wire2(100, 30)    <= sub_wire157(30);
	sub_wire2(100, 31)    <= sub_wire157(31);
	sub_wire2(100, 32)    <= sub_wire157(32);
	sub_wire2(100, 33)    <= sub_wire157(33);
	sub_wire2(100, 34)    <= sub_wire157(34);
	sub_wire2(100, 35)    <= sub_wire157(35);
	sub_wire2(100, 36)    <= sub_wire157(36);
	sub_wire2(100, 37)    <= sub_wire157(37);
	sub_wire2(100, 38)    <= sub_wire157(38);
	sub_wire2(100, 39)    <= sub_wire157(39);
	sub_wire2(99, 0)    <= sub_wire158(0);
	sub_wire2(99, 1)    <= sub_wire158(1);
	sub_wire2(99, 2)    <= sub_wire158(2);
	sub_wire2(99, 3)    <= sub_wire158(3);
	sub_wire2(99, 4)    <= sub_wire158(4);
	sub_wire2(99, 5)    <= sub_wire158(5);
	sub_wire2(99, 6)    <= sub_wire158(6);
	sub_wire2(99, 7)    <= sub_wire158(7);
	sub_wire2(99, 8)    <= sub_wire158(8);
	sub_wire2(99, 9)    <= sub_wire158(9);
	sub_wire2(99, 10)    <= sub_wire158(10);
	sub_wire2(99, 11)    <= sub_wire158(11);
	sub_wire2(99, 12)    <= sub_wire158(12);
	sub_wire2(99, 13)    <= sub_wire158(13);
	sub_wire2(99, 14)    <= sub_wire158(14);
	sub_wire2(99, 15)    <= sub_wire158(15);
	sub_wire2(99, 16)    <= sub_wire158(16);
	sub_wire2(99, 17)    <= sub_wire158(17);
	sub_wire2(99, 18)    <= sub_wire158(18);
	sub_wire2(99, 19)    <= sub_wire158(19);
	sub_wire2(99, 20)    <= sub_wire158(20);
	sub_wire2(99, 21)    <= sub_wire158(21);
	sub_wire2(99, 22)    <= sub_wire158(22);
	sub_wire2(99, 23)    <= sub_wire158(23);
	sub_wire2(99, 24)    <= sub_wire158(24);
	sub_wire2(99, 25)    <= sub_wire158(25);
	sub_wire2(99, 26)    <= sub_wire158(26);
	sub_wire2(99, 27)    <= sub_wire158(27);
	sub_wire2(99, 28)    <= sub_wire158(28);
	sub_wire2(99, 29)    <= sub_wire158(29);
	sub_wire2(99, 30)    <= sub_wire158(30);
	sub_wire2(99, 31)    <= sub_wire158(31);
	sub_wire2(99, 32)    <= sub_wire158(32);
	sub_wire2(99, 33)    <= sub_wire158(33);
	sub_wire2(99, 34)    <= sub_wire158(34);
	sub_wire2(99, 35)    <= sub_wire158(35);
	sub_wire2(99, 36)    <= sub_wire158(36);
	sub_wire2(99, 37)    <= sub_wire158(37);
	sub_wire2(99, 38)    <= sub_wire158(38);
	sub_wire2(99, 39)    <= sub_wire158(39);
	sub_wire2(98, 0)    <= sub_wire159(0);
	sub_wire2(98, 1)    <= sub_wire159(1);
	sub_wire2(98, 2)    <= sub_wire159(2);
	sub_wire2(98, 3)    <= sub_wire159(3);
	sub_wire2(98, 4)    <= sub_wire159(4);
	sub_wire2(98, 5)    <= sub_wire159(5);
	sub_wire2(98, 6)    <= sub_wire159(6);
	sub_wire2(98, 7)    <= sub_wire159(7);
	sub_wire2(98, 8)    <= sub_wire159(8);
	sub_wire2(98, 9)    <= sub_wire159(9);
	sub_wire2(98, 10)    <= sub_wire159(10);
	sub_wire2(98, 11)    <= sub_wire159(11);
	sub_wire2(98, 12)    <= sub_wire159(12);
	sub_wire2(98, 13)    <= sub_wire159(13);
	sub_wire2(98, 14)    <= sub_wire159(14);
	sub_wire2(98, 15)    <= sub_wire159(15);
	sub_wire2(98, 16)    <= sub_wire159(16);
	sub_wire2(98, 17)    <= sub_wire159(17);
	sub_wire2(98, 18)    <= sub_wire159(18);
	sub_wire2(98, 19)    <= sub_wire159(19);
	sub_wire2(98, 20)    <= sub_wire159(20);
	sub_wire2(98, 21)    <= sub_wire159(21);
	sub_wire2(98, 22)    <= sub_wire159(22);
	sub_wire2(98, 23)    <= sub_wire159(23);
	sub_wire2(98, 24)    <= sub_wire159(24);
	sub_wire2(98, 25)    <= sub_wire159(25);
	sub_wire2(98, 26)    <= sub_wire159(26);
	sub_wire2(98, 27)    <= sub_wire159(27);
	sub_wire2(98, 28)    <= sub_wire159(28);
	sub_wire2(98, 29)    <= sub_wire159(29);
	sub_wire2(98, 30)    <= sub_wire159(30);
	sub_wire2(98, 31)    <= sub_wire159(31);
	sub_wire2(98, 32)    <= sub_wire159(32);
	sub_wire2(98, 33)    <= sub_wire159(33);
	sub_wire2(98, 34)    <= sub_wire159(34);
	sub_wire2(98, 35)    <= sub_wire159(35);
	sub_wire2(98, 36)    <= sub_wire159(36);
	sub_wire2(98, 37)    <= sub_wire159(37);
	sub_wire2(98, 38)    <= sub_wire159(38);
	sub_wire2(98, 39)    <= sub_wire159(39);
	sub_wire2(97, 0)    <= sub_wire160(0);
	sub_wire2(97, 1)    <= sub_wire160(1);
	sub_wire2(97, 2)    <= sub_wire160(2);
	sub_wire2(97, 3)    <= sub_wire160(3);
	sub_wire2(97, 4)    <= sub_wire160(4);
	sub_wire2(97, 5)    <= sub_wire160(5);
	sub_wire2(97, 6)    <= sub_wire160(6);
	sub_wire2(97, 7)    <= sub_wire160(7);
	sub_wire2(97, 8)    <= sub_wire160(8);
	sub_wire2(97, 9)    <= sub_wire160(9);
	sub_wire2(97, 10)    <= sub_wire160(10);
	sub_wire2(97, 11)    <= sub_wire160(11);
	sub_wire2(97, 12)    <= sub_wire160(12);
	sub_wire2(97, 13)    <= sub_wire160(13);
	sub_wire2(97, 14)    <= sub_wire160(14);
	sub_wire2(97, 15)    <= sub_wire160(15);
	sub_wire2(97, 16)    <= sub_wire160(16);
	sub_wire2(97, 17)    <= sub_wire160(17);
	sub_wire2(97, 18)    <= sub_wire160(18);
	sub_wire2(97, 19)    <= sub_wire160(19);
	sub_wire2(97, 20)    <= sub_wire160(20);
	sub_wire2(97, 21)    <= sub_wire160(21);
	sub_wire2(97, 22)    <= sub_wire160(22);
	sub_wire2(97, 23)    <= sub_wire160(23);
	sub_wire2(97, 24)    <= sub_wire160(24);
	sub_wire2(97, 25)    <= sub_wire160(25);
	sub_wire2(97, 26)    <= sub_wire160(26);
	sub_wire2(97, 27)    <= sub_wire160(27);
	sub_wire2(97, 28)    <= sub_wire160(28);
	sub_wire2(97, 29)    <= sub_wire160(29);
	sub_wire2(97, 30)    <= sub_wire160(30);
	sub_wire2(97, 31)    <= sub_wire160(31);
	sub_wire2(97, 32)    <= sub_wire160(32);
	sub_wire2(97, 33)    <= sub_wire160(33);
	sub_wire2(97, 34)    <= sub_wire160(34);
	sub_wire2(97, 35)    <= sub_wire160(35);
	sub_wire2(97, 36)    <= sub_wire160(36);
	sub_wire2(97, 37)    <= sub_wire160(37);
	sub_wire2(97, 38)    <= sub_wire160(38);
	sub_wire2(97, 39)    <= sub_wire160(39);
	sub_wire2(96, 0)    <= sub_wire161(0);
	sub_wire2(96, 1)    <= sub_wire161(1);
	sub_wire2(96, 2)    <= sub_wire161(2);
	sub_wire2(96, 3)    <= sub_wire161(3);
	sub_wire2(96, 4)    <= sub_wire161(4);
	sub_wire2(96, 5)    <= sub_wire161(5);
	sub_wire2(96, 6)    <= sub_wire161(6);
	sub_wire2(96, 7)    <= sub_wire161(7);
	sub_wire2(96, 8)    <= sub_wire161(8);
	sub_wire2(96, 9)    <= sub_wire161(9);
	sub_wire2(96, 10)    <= sub_wire161(10);
	sub_wire2(96, 11)    <= sub_wire161(11);
	sub_wire2(96, 12)    <= sub_wire161(12);
	sub_wire2(96, 13)    <= sub_wire161(13);
	sub_wire2(96, 14)    <= sub_wire161(14);
	sub_wire2(96, 15)    <= sub_wire161(15);
	sub_wire2(96, 16)    <= sub_wire161(16);
	sub_wire2(96, 17)    <= sub_wire161(17);
	sub_wire2(96, 18)    <= sub_wire161(18);
	sub_wire2(96, 19)    <= sub_wire161(19);
	sub_wire2(96, 20)    <= sub_wire161(20);
	sub_wire2(96, 21)    <= sub_wire161(21);
	sub_wire2(96, 22)    <= sub_wire161(22);
	sub_wire2(96, 23)    <= sub_wire161(23);
	sub_wire2(96, 24)    <= sub_wire161(24);
	sub_wire2(96, 25)    <= sub_wire161(25);
	sub_wire2(96, 26)    <= sub_wire161(26);
	sub_wire2(96, 27)    <= sub_wire161(27);
	sub_wire2(96, 28)    <= sub_wire161(28);
	sub_wire2(96, 29)    <= sub_wire161(29);
	sub_wire2(96, 30)    <= sub_wire161(30);
	sub_wire2(96, 31)    <= sub_wire161(31);
	sub_wire2(96, 32)    <= sub_wire161(32);
	sub_wire2(96, 33)    <= sub_wire161(33);
	sub_wire2(96, 34)    <= sub_wire161(34);
	sub_wire2(96, 35)    <= sub_wire161(35);
	sub_wire2(96, 36)    <= sub_wire161(36);
	sub_wire2(96, 37)    <= sub_wire161(37);
	sub_wire2(96, 38)    <= sub_wire161(38);
	sub_wire2(96, 39)    <= sub_wire161(39);
	sub_wire2(95, 0)    <= sub_wire162(0);
	sub_wire2(95, 1)    <= sub_wire162(1);
	sub_wire2(95, 2)    <= sub_wire162(2);
	sub_wire2(95, 3)    <= sub_wire162(3);
	sub_wire2(95, 4)    <= sub_wire162(4);
	sub_wire2(95, 5)    <= sub_wire162(5);
	sub_wire2(95, 6)    <= sub_wire162(6);
	sub_wire2(95, 7)    <= sub_wire162(7);
	sub_wire2(95, 8)    <= sub_wire162(8);
	sub_wire2(95, 9)    <= sub_wire162(9);
	sub_wire2(95, 10)    <= sub_wire162(10);
	sub_wire2(95, 11)    <= sub_wire162(11);
	sub_wire2(95, 12)    <= sub_wire162(12);
	sub_wire2(95, 13)    <= sub_wire162(13);
	sub_wire2(95, 14)    <= sub_wire162(14);
	sub_wire2(95, 15)    <= sub_wire162(15);
	sub_wire2(95, 16)    <= sub_wire162(16);
	sub_wire2(95, 17)    <= sub_wire162(17);
	sub_wire2(95, 18)    <= sub_wire162(18);
	sub_wire2(95, 19)    <= sub_wire162(19);
	sub_wire2(95, 20)    <= sub_wire162(20);
	sub_wire2(95, 21)    <= sub_wire162(21);
	sub_wire2(95, 22)    <= sub_wire162(22);
	sub_wire2(95, 23)    <= sub_wire162(23);
	sub_wire2(95, 24)    <= sub_wire162(24);
	sub_wire2(95, 25)    <= sub_wire162(25);
	sub_wire2(95, 26)    <= sub_wire162(26);
	sub_wire2(95, 27)    <= sub_wire162(27);
	sub_wire2(95, 28)    <= sub_wire162(28);
	sub_wire2(95, 29)    <= sub_wire162(29);
	sub_wire2(95, 30)    <= sub_wire162(30);
	sub_wire2(95, 31)    <= sub_wire162(31);
	sub_wire2(95, 32)    <= sub_wire162(32);
	sub_wire2(95, 33)    <= sub_wire162(33);
	sub_wire2(95, 34)    <= sub_wire162(34);
	sub_wire2(95, 35)    <= sub_wire162(35);
	sub_wire2(95, 36)    <= sub_wire162(36);
	sub_wire2(95, 37)    <= sub_wire162(37);
	sub_wire2(95, 38)    <= sub_wire162(38);
	sub_wire2(95, 39)    <= sub_wire162(39);
	sub_wire2(94, 0)    <= sub_wire163(0);
	sub_wire2(94, 1)    <= sub_wire163(1);
	sub_wire2(94, 2)    <= sub_wire163(2);
	sub_wire2(94, 3)    <= sub_wire163(3);
	sub_wire2(94, 4)    <= sub_wire163(4);
	sub_wire2(94, 5)    <= sub_wire163(5);
	sub_wire2(94, 6)    <= sub_wire163(6);
	sub_wire2(94, 7)    <= sub_wire163(7);
	sub_wire2(94, 8)    <= sub_wire163(8);
	sub_wire2(94, 9)    <= sub_wire163(9);
	sub_wire2(94, 10)    <= sub_wire163(10);
	sub_wire2(94, 11)    <= sub_wire163(11);
	sub_wire2(94, 12)    <= sub_wire163(12);
	sub_wire2(94, 13)    <= sub_wire163(13);
	sub_wire2(94, 14)    <= sub_wire163(14);
	sub_wire2(94, 15)    <= sub_wire163(15);
	sub_wire2(94, 16)    <= sub_wire163(16);
	sub_wire2(94, 17)    <= sub_wire163(17);
	sub_wire2(94, 18)    <= sub_wire163(18);
	sub_wire2(94, 19)    <= sub_wire163(19);
	sub_wire2(94, 20)    <= sub_wire163(20);
	sub_wire2(94, 21)    <= sub_wire163(21);
	sub_wire2(94, 22)    <= sub_wire163(22);
	sub_wire2(94, 23)    <= sub_wire163(23);
	sub_wire2(94, 24)    <= sub_wire163(24);
	sub_wire2(94, 25)    <= sub_wire163(25);
	sub_wire2(94, 26)    <= sub_wire163(26);
	sub_wire2(94, 27)    <= sub_wire163(27);
	sub_wire2(94, 28)    <= sub_wire163(28);
	sub_wire2(94, 29)    <= sub_wire163(29);
	sub_wire2(94, 30)    <= sub_wire163(30);
	sub_wire2(94, 31)    <= sub_wire163(31);
	sub_wire2(94, 32)    <= sub_wire163(32);
	sub_wire2(94, 33)    <= sub_wire163(33);
	sub_wire2(94, 34)    <= sub_wire163(34);
	sub_wire2(94, 35)    <= sub_wire163(35);
	sub_wire2(94, 36)    <= sub_wire163(36);
	sub_wire2(94, 37)    <= sub_wire163(37);
	sub_wire2(94, 38)    <= sub_wire163(38);
	sub_wire2(94, 39)    <= sub_wire163(39);
	sub_wire2(93, 0)    <= sub_wire164(0);
	sub_wire2(93, 1)    <= sub_wire164(1);
	sub_wire2(93, 2)    <= sub_wire164(2);
	sub_wire2(93, 3)    <= sub_wire164(3);
	sub_wire2(93, 4)    <= sub_wire164(4);
	sub_wire2(93, 5)    <= sub_wire164(5);
	sub_wire2(93, 6)    <= sub_wire164(6);
	sub_wire2(93, 7)    <= sub_wire164(7);
	sub_wire2(93, 8)    <= sub_wire164(8);
	sub_wire2(93, 9)    <= sub_wire164(9);
	sub_wire2(93, 10)    <= sub_wire164(10);
	sub_wire2(93, 11)    <= sub_wire164(11);
	sub_wire2(93, 12)    <= sub_wire164(12);
	sub_wire2(93, 13)    <= sub_wire164(13);
	sub_wire2(93, 14)    <= sub_wire164(14);
	sub_wire2(93, 15)    <= sub_wire164(15);
	sub_wire2(93, 16)    <= sub_wire164(16);
	sub_wire2(93, 17)    <= sub_wire164(17);
	sub_wire2(93, 18)    <= sub_wire164(18);
	sub_wire2(93, 19)    <= sub_wire164(19);
	sub_wire2(93, 20)    <= sub_wire164(20);
	sub_wire2(93, 21)    <= sub_wire164(21);
	sub_wire2(93, 22)    <= sub_wire164(22);
	sub_wire2(93, 23)    <= sub_wire164(23);
	sub_wire2(93, 24)    <= sub_wire164(24);
	sub_wire2(93, 25)    <= sub_wire164(25);
	sub_wire2(93, 26)    <= sub_wire164(26);
	sub_wire2(93, 27)    <= sub_wire164(27);
	sub_wire2(93, 28)    <= sub_wire164(28);
	sub_wire2(93, 29)    <= sub_wire164(29);
	sub_wire2(93, 30)    <= sub_wire164(30);
	sub_wire2(93, 31)    <= sub_wire164(31);
	sub_wire2(93, 32)    <= sub_wire164(32);
	sub_wire2(93, 33)    <= sub_wire164(33);
	sub_wire2(93, 34)    <= sub_wire164(34);
	sub_wire2(93, 35)    <= sub_wire164(35);
	sub_wire2(93, 36)    <= sub_wire164(36);
	sub_wire2(93, 37)    <= sub_wire164(37);
	sub_wire2(93, 38)    <= sub_wire164(38);
	sub_wire2(93, 39)    <= sub_wire164(39);
	sub_wire2(92, 0)    <= sub_wire165(0);
	sub_wire2(92, 1)    <= sub_wire165(1);
	sub_wire2(92, 2)    <= sub_wire165(2);
	sub_wire2(92, 3)    <= sub_wire165(3);
	sub_wire2(92, 4)    <= sub_wire165(4);
	sub_wire2(92, 5)    <= sub_wire165(5);
	sub_wire2(92, 6)    <= sub_wire165(6);
	sub_wire2(92, 7)    <= sub_wire165(7);
	sub_wire2(92, 8)    <= sub_wire165(8);
	sub_wire2(92, 9)    <= sub_wire165(9);
	sub_wire2(92, 10)    <= sub_wire165(10);
	sub_wire2(92, 11)    <= sub_wire165(11);
	sub_wire2(92, 12)    <= sub_wire165(12);
	sub_wire2(92, 13)    <= sub_wire165(13);
	sub_wire2(92, 14)    <= sub_wire165(14);
	sub_wire2(92, 15)    <= sub_wire165(15);
	sub_wire2(92, 16)    <= sub_wire165(16);
	sub_wire2(92, 17)    <= sub_wire165(17);
	sub_wire2(92, 18)    <= sub_wire165(18);
	sub_wire2(92, 19)    <= sub_wire165(19);
	sub_wire2(92, 20)    <= sub_wire165(20);
	sub_wire2(92, 21)    <= sub_wire165(21);
	sub_wire2(92, 22)    <= sub_wire165(22);
	sub_wire2(92, 23)    <= sub_wire165(23);
	sub_wire2(92, 24)    <= sub_wire165(24);
	sub_wire2(92, 25)    <= sub_wire165(25);
	sub_wire2(92, 26)    <= sub_wire165(26);
	sub_wire2(92, 27)    <= sub_wire165(27);
	sub_wire2(92, 28)    <= sub_wire165(28);
	sub_wire2(92, 29)    <= sub_wire165(29);
	sub_wire2(92, 30)    <= sub_wire165(30);
	sub_wire2(92, 31)    <= sub_wire165(31);
	sub_wire2(92, 32)    <= sub_wire165(32);
	sub_wire2(92, 33)    <= sub_wire165(33);
	sub_wire2(92, 34)    <= sub_wire165(34);
	sub_wire2(92, 35)    <= sub_wire165(35);
	sub_wire2(92, 36)    <= sub_wire165(36);
	sub_wire2(92, 37)    <= sub_wire165(37);
	sub_wire2(92, 38)    <= sub_wire165(38);
	sub_wire2(92, 39)    <= sub_wire165(39);
	sub_wire2(91, 0)    <= sub_wire166(0);
	sub_wire2(91, 1)    <= sub_wire166(1);
	sub_wire2(91, 2)    <= sub_wire166(2);
	sub_wire2(91, 3)    <= sub_wire166(3);
	sub_wire2(91, 4)    <= sub_wire166(4);
	sub_wire2(91, 5)    <= sub_wire166(5);
	sub_wire2(91, 6)    <= sub_wire166(6);
	sub_wire2(91, 7)    <= sub_wire166(7);
	sub_wire2(91, 8)    <= sub_wire166(8);
	sub_wire2(91, 9)    <= sub_wire166(9);
	sub_wire2(91, 10)    <= sub_wire166(10);
	sub_wire2(91, 11)    <= sub_wire166(11);
	sub_wire2(91, 12)    <= sub_wire166(12);
	sub_wire2(91, 13)    <= sub_wire166(13);
	sub_wire2(91, 14)    <= sub_wire166(14);
	sub_wire2(91, 15)    <= sub_wire166(15);
	sub_wire2(91, 16)    <= sub_wire166(16);
	sub_wire2(91, 17)    <= sub_wire166(17);
	sub_wire2(91, 18)    <= sub_wire166(18);
	sub_wire2(91, 19)    <= sub_wire166(19);
	sub_wire2(91, 20)    <= sub_wire166(20);
	sub_wire2(91, 21)    <= sub_wire166(21);
	sub_wire2(91, 22)    <= sub_wire166(22);
	sub_wire2(91, 23)    <= sub_wire166(23);
	sub_wire2(91, 24)    <= sub_wire166(24);
	sub_wire2(91, 25)    <= sub_wire166(25);
	sub_wire2(91, 26)    <= sub_wire166(26);
	sub_wire2(91, 27)    <= sub_wire166(27);
	sub_wire2(91, 28)    <= sub_wire166(28);
	sub_wire2(91, 29)    <= sub_wire166(29);
	sub_wire2(91, 30)    <= sub_wire166(30);
	sub_wire2(91, 31)    <= sub_wire166(31);
	sub_wire2(91, 32)    <= sub_wire166(32);
	sub_wire2(91, 33)    <= sub_wire166(33);
	sub_wire2(91, 34)    <= sub_wire166(34);
	sub_wire2(91, 35)    <= sub_wire166(35);
	sub_wire2(91, 36)    <= sub_wire166(36);
	sub_wire2(91, 37)    <= sub_wire166(37);
	sub_wire2(91, 38)    <= sub_wire166(38);
	sub_wire2(91, 39)    <= sub_wire166(39);
	sub_wire2(90, 0)    <= sub_wire167(0);
	sub_wire2(90, 1)    <= sub_wire167(1);
	sub_wire2(90, 2)    <= sub_wire167(2);
	sub_wire2(90, 3)    <= sub_wire167(3);
	sub_wire2(90, 4)    <= sub_wire167(4);
	sub_wire2(90, 5)    <= sub_wire167(5);
	sub_wire2(90, 6)    <= sub_wire167(6);
	sub_wire2(90, 7)    <= sub_wire167(7);
	sub_wire2(90, 8)    <= sub_wire167(8);
	sub_wire2(90, 9)    <= sub_wire167(9);
	sub_wire2(90, 10)    <= sub_wire167(10);
	sub_wire2(90, 11)    <= sub_wire167(11);
	sub_wire2(90, 12)    <= sub_wire167(12);
	sub_wire2(90, 13)    <= sub_wire167(13);
	sub_wire2(90, 14)    <= sub_wire167(14);
	sub_wire2(90, 15)    <= sub_wire167(15);
	sub_wire2(90, 16)    <= sub_wire167(16);
	sub_wire2(90, 17)    <= sub_wire167(17);
	sub_wire2(90, 18)    <= sub_wire167(18);
	sub_wire2(90, 19)    <= sub_wire167(19);
	sub_wire2(90, 20)    <= sub_wire167(20);
	sub_wire2(90, 21)    <= sub_wire167(21);
	sub_wire2(90, 22)    <= sub_wire167(22);
	sub_wire2(90, 23)    <= sub_wire167(23);
	sub_wire2(90, 24)    <= sub_wire167(24);
	sub_wire2(90, 25)    <= sub_wire167(25);
	sub_wire2(90, 26)    <= sub_wire167(26);
	sub_wire2(90, 27)    <= sub_wire167(27);
	sub_wire2(90, 28)    <= sub_wire167(28);
	sub_wire2(90, 29)    <= sub_wire167(29);
	sub_wire2(90, 30)    <= sub_wire167(30);
	sub_wire2(90, 31)    <= sub_wire167(31);
	sub_wire2(90, 32)    <= sub_wire167(32);
	sub_wire2(90, 33)    <= sub_wire167(33);
	sub_wire2(90, 34)    <= sub_wire167(34);
	sub_wire2(90, 35)    <= sub_wire167(35);
	sub_wire2(90, 36)    <= sub_wire167(36);
	sub_wire2(90, 37)    <= sub_wire167(37);
	sub_wire2(90, 38)    <= sub_wire167(38);
	sub_wire2(90, 39)    <= sub_wire167(39);
	sub_wire2(89, 0)    <= sub_wire168(0);
	sub_wire2(89, 1)    <= sub_wire168(1);
	sub_wire2(89, 2)    <= sub_wire168(2);
	sub_wire2(89, 3)    <= sub_wire168(3);
	sub_wire2(89, 4)    <= sub_wire168(4);
	sub_wire2(89, 5)    <= sub_wire168(5);
	sub_wire2(89, 6)    <= sub_wire168(6);
	sub_wire2(89, 7)    <= sub_wire168(7);
	sub_wire2(89, 8)    <= sub_wire168(8);
	sub_wire2(89, 9)    <= sub_wire168(9);
	sub_wire2(89, 10)    <= sub_wire168(10);
	sub_wire2(89, 11)    <= sub_wire168(11);
	sub_wire2(89, 12)    <= sub_wire168(12);
	sub_wire2(89, 13)    <= sub_wire168(13);
	sub_wire2(89, 14)    <= sub_wire168(14);
	sub_wire2(89, 15)    <= sub_wire168(15);
	sub_wire2(89, 16)    <= sub_wire168(16);
	sub_wire2(89, 17)    <= sub_wire168(17);
	sub_wire2(89, 18)    <= sub_wire168(18);
	sub_wire2(89, 19)    <= sub_wire168(19);
	sub_wire2(89, 20)    <= sub_wire168(20);
	sub_wire2(89, 21)    <= sub_wire168(21);
	sub_wire2(89, 22)    <= sub_wire168(22);
	sub_wire2(89, 23)    <= sub_wire168(23);
	sub_wire2(89, 24)    <= sub_wire168(24);
	sub_wire2(89, 25)    <= sub_wire168(25);
	sub_wire2(89, 26)    <= sub_wire168(26);
	sub_wire2(89, 27)    <= sub_wire168(27);
	sub_wire2(89, 28)    <= sub_wire168(28);
	sub_wire2(89, 29)    <= sub_wire168(29);
	sub_wire2(89, 30)    <= sub_wire168(30);
	sub_wire2(89, 31)    <= sub_wire168(31);
	sub_wire2(89, 32)    <= sub_wire168(32);
	sub_wire2(89, 33)    <= sub_wire168(33);
	sub_wire2(89, 34)    <= sub_wire168(34);
	sub_wire2(89, 35)    <= sub_wire168(35);
	sub_wire2(89, 36)    <= sub_wire168(36);
	sub_wire2(89, 37)    <= sub_wire168(37);
	sub_wire2(89, 38)    <= sub_wire168(38);
	sub_wire2(89, 39)    <= sub_wire168(39);
	sub_wire2(88, 0)    <= sub_wire169(0);
	sub_wire2(88, 1)    <= sub_wire169(1);
	sub_wire2(88, 2)    <= sub_wire169(2);
	sub_wire2(88, 3)    <= sub_wire169(3);
	sub_wire2(88, 4)    <= sub_wire169(4);
	sub_wire2(88, 5)    <= sub_wire169(5);
	sub_wire2(88, 6)    <= sub_wire169(6);
	sub_wire2(88, 7)    <= sub_wire169(7);
	sub_wire2(88, 8)    <= sub_wire169(8);
	sub_wire2(88, 9)    <= sub_wire169(9);
	sub_wire2(88, 10)    <= sub_wire169(10);
	sub_wire2(88, 11)    <= sub_wire169(11);
	sub_wire2(88, 12)    <= sub_wire169(12);
	sub_wire2(88, 13)    <= sub_wire169(13);
	sub_wire2(88, 14)    <= sub_wire169(14);
	sub_wire2(88, 15)    <= sub_wire169(15);
	sub_wire2(88, 16)    <= sub_wire169(16);
	sub_wire2(88, 17)    <= sub_wire169(17);
	sub_wire2(88, 18)    <= sub_wire169(18);
	sub_wire2(88, 19)    <= sub_wire169(19);
	sub_wire2(88, 20)    <= sub_wire169(20);
	sub_wire2(88, 21)    <= sub_wire169(21);
	sub_wire2(88, 22)    <= sub_wire169(22);
	sub_wire2(88, 23)    <= sub_wire169(23);
	sub_wire2(88, 24)    <= sub_wire169(24);
	sub_wire2(88, 25)    <= sub_wire169(25);
	sub_wire2(88, 26)    <= sub_wire169(26);
	sub_wire2(88, 27)    <= sub_wire169(27);
	sub_wire2(88, 28)    <= sub_wire169(28);
	sub_wire2(88, 29)    <= sub_wire169(29);
	sub_wire2(88, 30)    <= sub_wire169(30);
	sub_wire2(88, 31)    <= sub_wire169(31);
	sub_wire2(88, 32)    <= sub_wire169(32);
	sub_wire2(88, 33)    <= sub_wire169(33);
	sub_wire2(88, 34)    <= sub_wire169(34);
	sub_wire2(88, 35)    <= sub_wire169(35);
	sub_wire2(88, 36)    <= sub_wire169(36);
	sub_wire2(88, 37)    <= sub_wire169(37);
	sub_wire2(88, 38)    <= sub_wire169(38);
	sub_wire2(88, 39)    <= sub_wire169(39);
	sub_wire2(87, 0)    <= sub_wire170(0);
	sub_wire2(87, 1)    <= sub_wire170(1);
	sub_wire2(87, 2)    <= sub_wire170(2);
	sub_wire2(87, 3)    <= sub_wire170(3);
	sub_wire2(87, 4)    <= sub_wire170(4);
	sub_wire2(87, 5)    <= sub_wire170(5);
	sub_wire2(87, 6)    <= sub_wire170(6);
	sub_wire2(87, 7)    <= sub_wire170(7);
	sub_wire2(87, 8)    <= sub_wire170(8);
	sub_wire2(87, 9)    <= sub_wire170(9);
	sub_wire2(87, 10)    <= sub_wire170(10);
	sub_wire2(87, 11)    <= sub_wire170(11);
	sub_wire2(87, 12)    <= sub_wire170(12);
	sub_wire2(87, 13)    <= sub_wire170(13);
	sub_wire2(87, 14)    <= sub_wire170(14);
	sub_wire2(87, 15)    <= sub_wire170(15);
	sub_wire2(87, 16)    <= sub_wire170(16);
	sub_wire2(87, 17)    <= sub_wire170(17);
	sub_wire2(87, 18)    <= sub_wire170(18);
	sub_wire2(87, 19)    <= sub_wire170(19);
	sub_wire2(87, 20)    <= sub_wire170(20);
	sub_wire2(87, 21)    <= sub_wire170(21);
	sub_wire2(87, 22)    <= sub_wire170(22);
	sub_wire2(87, 23)    <= sub_wire170(23);
	sub_wire2(87, 24)    <= sub_wire170(24);
	sub_wire2(87, 25)    <= sub_wire170(25);
	sub_wire2(87, 26)    <= sub_wire170(26);
	sub_wire2(87, 27)    <= sub_wire170(27);
	sub_wire2(87, 28)    <= sub_wire170(28);
	sub_wire2(87, 29)    <= sub_wire170(29);
	sub_wire2(87, 30)    <= sub_wire170(30);
	sub_wire2(87, 31)    <= sub_wire170(31);
	sub_wire2(87, 32)    <= sub_wire170(32);
	sub_wire2(87, 33)    <= sub_wire170(33);
	sub_wire2(87, 34)    <= sub_wire170(34);
	sub_wire2(87, 35)    <= sub_wire170(35);
	sub_wire2(87, 36)    <= sub_wire170(36);
	sub_wire2(87, 37)    <= sub_wire170(37);
	sub_wire2(87, 38)    <= sub_wire170(38);
	sub_wire2(87, 39)    <= sub_wire170(39);
	sub_wire2(86, 0)    <= sub_wire171(0);
	sub_wire2(86, 1)    <= sub_wire171(1);
	sub_wire2(86, 2)    <= sub_wire171(2);
	sub_wire2(86, 3)    <= sub_wire171(3);
	sub_wire2(86, 4)    <= sub_wire171(4);
	sub_wire2(86, 5)    <= sub_wire171(5);
	sub_wire2(86, 6)    <= sub_wire171(6);
	sub_wire2(86, 7)    <= sub_wire171(7);
	sub_wire2(86, 8)    <= sub_wire171(8);
	sub_wire2(86, 9)    <= sub_wire171(9);
	sub_wire2(86, 10)    <= sub_wire171(10);
	sub_wire2(86, 11)    <= sub_wire171(11);
	sub_wire2(86, 12)    <= sub_wire171(12);
	sub_wire2(86, 13)    <= sub_wire171(13);
	sub_wire2(86, 14)    <= sub_wire171(14);
	sub_wire2(86, 15)    <= sub_wire171(15);
	sub_wire2(86, 16)    <= sub_wire171(16);
	sub_wire2(86, 17)    <= sub_wire171(17);
	sub_wire2(86, 18)    <= sub_wire171(18);
	sub_wire2(86, 19)    <= sub_wire171(19);
	sub_wire2(86, 20)    <= sub_wire171(20);
	sub_wire2(86, 21)    <= sub_wire171(21);
	sub_wire2(86, 22)    <= sub_wire171(22);
	sub_wire2(86, 23)    <= sub_wire171(23);
	sub_wire2(86, 24)    <= sub_wire171(24);
	sub_wire2(86, 25)    <= sub_wire171(25);
	sub_wire2(86, 26)    <= sub_wire171(26);
	sub_wire2(86, 27)    <= sub_wire171(27);
	sub_wire2(86, 28)    <= sub_wire171(28);
	sub_wire2(86, 29)    <= sub_wire171(29);
	sub_wire2(86, 30)    <= sub_wire171(30);
	sub_wire2(86, 31)    <= sub_wire171(31);
	sub_wire2(86, 32)    <= sub_wire171(32);
	sub_wire2(86, 33)    <= sub_wire171(33);
	sub_wire2(86, 34)    <= sub_wire171(34);
	sub_wire2(86, 35)    <= sub_wire171(35);
	sub_wire2(86, 36)    <= sub_wire171(36);
	sub_wire2(86, 37)    <= sub_wire171(37);
	sub_wire2(86, 38)    <= sub_wire171(38);
	sub_wire2(86, 39)    <= sub_wire171(39);
	sub_wire2(85, 0)    <= sub_wire172(0);
	sub_wire2(85, 1)    <= sub_wire172(1);
	sub_wire2(85, 2)    <= sub_wire172(2);
	sub_wire2(85, 3)    <= sub_wire172(3);
	sub_wire2(85, 4)    <= sub_wire172(4);
	sub_wire2(85, 5)    <= sub_wire172(5);
	sub_wire2(85, 6)    <= sub_wire172(6);
	sub_wire2(85, 7)    <= sub_wire172(7);
	sub_wire2(85, 8)    <= sub_wire172(8);
	sub_wire2(85, 9)    <= sub_wire172(9);
	sub_wire2(85, 10)    <= sub_wire172(10);
	sub_wire2(85, 11)    <= sub_wire172(11);
	sub_wire2(85, 12)    <= sub_wire172(12);
	sub_wire2(85, 13)    <= sub_wire172(13);
	sub_wire2(85, 14)    <= sub_wire172(14);
	sub_wire2(85, 15)    <= sub_wire172(15);
	sub_wire2(85, 16)    <= sub_wire172(16);
	sub_wire2(85, 17)    <= sub_wire172(17);
	sub_wire2(85, 18)    <= sub_wire172(18);
	sub_wire2(85, 19)    <= sub_wire172(19);
	sub_wire2(85, 20)    <= sub_wire172(20);
	sub_wire2(85, 21)    <= sub_wire172(21);
	sub_wire2(85, 22)    <= sub_wire172(22);
	sub_wire2(85, 23)    <= sub_wire172(23);
	sub_wire2(85, 24)    <= sub_wire172(24);
	sub_wire2(85, 25)    <= sub_wire172(25);
	sub_wire2(85, 26)    <= sub_wire172(26);
	sub_wire2(85, 27)    <= sub_wire172(27);
	sub_wire2(85, 28)    <= sub_wire172(28);
	sub_wire2(85, 29)    <= sub_wire172(29);
	sub_wire2(85, 30)    <= sub_wire172(30);
	sub_wire2(85, 31)    <= sub_wire172(31);
	sub_wire2(85, 32)    <= sub_wire172(32);
	sub_wire2(85, 33)    <= sub_wire172(33);
	sub_wire2(85, 34)    <= sub_wire172(34);
	sub_wire2(85, 35)    <= sub_wire172(35);
	sub_wire2(85, 36)    <= sub_wire172(36);
	sub_wire2(85, 37)    <= sub_wire172(37);
	sub_wire2(85, 38)    <= sub_wire172(38);
	sub_wire2(85, 39)    <= sub_wire172(39);
	sub_wire2(84, 0)    <= sub_wire173(0);
	sub_wire2(84, 1)    <= sub_wire173(1);
	sub_wire2(84, 2)    <= sub_wire173(2);
	sub_wire2(84, 3)    <= sub_wire173(3);
	sub_wire2(84, 4)    <= sub_wire173(4);
	sub_wire2(84, 5)    <= sub_wire173(5);
	sub_wire2(84, 6)    <= sub_wire173(6);
	sub_wire2(84, 7)    <= sub_wire173(7);
	sub_wire2(84, 8)    <= sub_wire173(8);
	sub_wire2(84, 9)    <= sub_wire173(9);
	sub_wire2(84, 10)    <= sub_wire173(10);
	sub_wire2(84, 11)    <= sub_wire173(11);
	sub_wire2(84, 12)    <= sub_wire173(12);
	sub_wire2(84, 13)    <= sub_wire173(13);
	sub_wire2(84, 14)    <= sub_wire173(14);
	sub_wire2(84, 15)    <= sub_wire173(15);
	sub_wire2(84, 16)    <= sub_wire173(16);
	sub_wire2(84, 17)    <= sub_wire173(17);
	sub_wire2(84, 18)    <= sub_wire173(18);
	sub_wire2(84, 19)    <= sub_wire173(19);
	sub_wire2(84, 20)    <= sub_wire173(20);
	sub_wire2(84, 21)    <= sub_wire173(21);
	sub_wire2(84, 22)    <= sub_wire173(22);
	sub_wire2(84, 23)    <= sub_wire173(23);
	sub_wire2(84, 24)    <= sub_wire173(24);
	sub_wire2(84, 25)    <= sub_wire173(25);
	sub_wire2(84, 26)    <= sub_wire173(26);
	sub_wire2(84, 27)    <= sub_wire173(27);
	sub_wire2(84, 28)    <= sub_wire173(28);
	sub_wire2(84, 29)    <= sub_wire173(29);
	sub_wire2(84, 30)    <= sub_wire173(30);
	sub_wire2(84, 31)    <= sub_wire173(31);
	sub_wire2(84, 32)    <= sub_wire173(32);
	sub_wire2(84, 33)    <= sub_wire173(33);
	sub_wire2(84, 34)    <= sub_wire173(34);
	sub_wire2(84, 35)    <= sub_wire173(35);
	sub_wire2(84, 36)    <= sub_wire173(36);
	sub_wire2(84, 37)    <= sub_wire173(37);
	sub_wire2(84, 38)    <= sub_wire173(38);
	sub_wire2(84, 39)    <= sub_wire173(39);
	sub_wire2(83, 0)    <= sub_wire174(0);
	sub_wire2(83, 1)    <= sub_wire174(1);
	sub_wire2(83, 2)    <= sub_wire174(2);
	sub_wire2(83, 3)    <= sub_wire174(3);
	sub_wire2(83, 4)    <= sub_wire174(4);
	sub_wire2(83, 5)    <= sub_wire174(5);
	sub_wire2(83, 6)    <= sub_wire174(6);
	sub_wire2(83, 7)    <= sub_wire174(7);
	sub_wire2(83, 8)    <= sub_wire174(8);
	sub_wire2(83, 9)    <= sub_wire174(9);
	sub_wire2(83, 10)    <= sub_wire174(10);
	sub_wire2(83, 11)    <= sub_wire174(11);
	sub_wire2(83, 12)    <= sub_wire174(12);
	sub_wire2(83, 13)    <= sub_wire174(13);
	sub_wire2(83, 14)    <= sub_wire174(14);
	sub_wire2(83, 15)    <= sub_wire174(15);
	sub_wire2(83, 16)    <= sub_wire174(16);
	sub_wire2(83, 17)    <= sub_wire174(17);
	sub_wire2(83, 18)    <= sub_wire174(18);
	sub_wire2(83, 19)    <= sub_wire174(19);
	sub_wire2(83, 20)    <= sub_wire174(20);
	sub_wire2(83, 21)    <= sub_wire174(21);
	sub_wire2(83, 22)    <= sub_wire174(22);
	sub_wire2(83, 23)    <= sub_wire174(23);
	sub_wire2(83, 24)    <= sub_wire174(24);
	sub_wire2(83, 25)    <= sub_wire174(25);
	sub_wire2(83, 26)    <= sub_wire174(26);
	sub_wire2(83, 27)    <= sub_wire174(27);
	sub_wire2(83, 28)    <= sub_wire174(28);
	sub_wire2(83, 29)    <= sub_wire174(29);
	sub_wire2(83, 30)    <= sub_wire174(30);
	sub_wire2(83, 31)    <= sub_wire174(31);
	sub_wire2(83, 32)    <= sub_wire174(32);
	sub_wire2(83, 33)    <= sub_wire174(33);
	sub_wire2(83, 34)    <= sub_wire174(34);
	sub_wire2(83, 35)    <= sub_wire174(35);
	sub_wire2(83, 36)    <= sub_wire174(36);
	sub_wire2(83, 37)    <= sub_wire174(37);
	sub_wire2(83, 38)    <= sub_wire174(38);
	sub_wire2(83, 39)    <= sub_wire174(39);
	sub_wire2(82, 0)    <= sub_wire175(0);
	sub_wire2(82, 1)    <= sub_wire175(1);
	sub_wire2(82, 2)    <= sub_wire175(2);
	sub_wire2(82, 3)    <= sub_wire175(3);
	sub_wire2(82, 4)    <= sub_wire175(4);
	sub_wire2(82, 5)    <= sub_wire175(5);
	sub_wire2(82, 6)    <= sub_wire175(6);
	sub_wire2(82, 7)    <= sub_wire175(7);
	sub_wire2(82, 8)    <= sub_wire175(8);
	sub_wire2(82, 9)    <= sub_wire175(9);
	sub_wire2(82, 10)    <= sub_wire175(10);
	sub_wire2(82, 11)    <= sub_wire175(11);
	sub_wire2(82, 12)    <= sub_wire175(12);
	sub_wire2(82, 13)    <= sub_wire175(13);
	sub_wire2(82, 14)    <= sub_wire175(14);
	sub_wire2(82, 15)    <= sub_wire175(15);
	sub_wire2(82, 16)    <= sub_wire175(16);
	sub_wire2(82, 17)    <= sub_wire175(17);
	sub_wire2(82, 18)    <= sub_wire175(18);
	sub_wire2(82, 19)    <= sub_wire175(19);
	sub_wire2(82, 20)    <= sub_wire175(20);
	sub_wire2(82, 21)    <= sub_wire175(21);
	sub_wire2(82, 22)    <= sub_wire175(22);
	sub_wire2(82, 23)    <= sub_wire175(23);
	sub_wire2(82, 24)    <= sub_wire175(24);
	sub_wire2(82, 25)    <= sub_wire175(25);
	sub_wire2(82, 26)    <= sub_wire175(26);
	sub_wire2(82, 27)    <= sub_wire175(27);
	sub_wire2(82, 28)    <= sub_wire175(28);
	sub_wire2(82, 29)    <= sub_wire175(29);
	sub_wire2(82, 30)    <= sub_wire175(30);
	sub_wire2(82, 31)    <= sub_wire175(31);
	sub_wire2(82, 32)    <= sub_wire175(32);
	sub_wire2(82, 33)    <= sub_wire175(33);
	sub_wire2(82, 34)    <= sub_wire175(34);
	sub_wire2(82, 35)    <= sub_wire175(35);
	sub_wire2(82, 36)    <= sub_wire175(36);
	sub_wire2(82, 37)    <= sub_wire175(37);
	sub_wire2(82, 38)    <= sub_wire175(38);
	sub_wire2(82, 39)    <= sub_wire175(39);
	sub_wire2(81, 0)    <= sub_wire176(0);
	sub_wire2(81, 1)    <= sub_wire176(1);
	sub_wire2(81, 2)    <= sub_wire176(2);
	sub_wire2(81, 3)    <= sub_wire176(3);
	sub_wire2(81, 4)    <= sub_wire176(4);
	sub_wire2(81, 5)    <= sub_wire176(5);
	sub_wire2(81, 6)    <= sub_wire176(6);
	sub_wire2(81, 7)    <= sub_wire176(7);
	sub_wire2(81, 8)    <= sub_wire176(8);
	sub_wire2(81, 9)    <= sub_wire176(9);
	sub_wire2(81, 10)    <= sub_wire176(10);
	sub_wire2(81, 11)    <= sub_wire176(11);
	sub_wire2(81, 12)    <= sub_wire176(12);
	sub_wire2(81, 13)    <= sub_wire176(13);
	sub_wire2(81, 14)    <= sub_wire176(14);
	sub_wire2(81, 15)    <= sub_wire176(15);
	sub_wire2(81, 16)    <= sub_wire176(16);
	sub_wire2(81, 17)    <= sub_wire176(17);
	sub_wire2(81, 18)    <= sub_wire176(18);
	sub_wire2(81, 19)    <= sub_wire176(19);
	sub_wire2(81, 20)    <= sub_wire176(20);
	sub_wire2(81, 21)    <= sub_wire176(21);
	sub_wire2(81, 22)    <= sub_wire176(22);
	sub_wire2(81, 23)    <= sub_wire176(23);
	sub_wire2(81, 24)    <= sub_wire176(24);
	sub_wire2(81, 25)    <= sub_wire176(25);
	sub_wire2(81, 26)    <= sub_wire176(26);
	sub_wire2(81, 27)    <= sub_wire176(27);
	sub_wire2(81, 28)    <= sub_wire176(28);
	sub_wire2(81, 29)    <= sub_wire176(29);
	sub_wire2(81, 30)    <= sub_wire176(30);
	sub_wire2(81, 31)    <= sub_wire176(31);
	sub_wire2(81, 32)    <= sub_wire176(32);
	sub_wire2(81, 33)    <= sub_wire176(33);
	sub_wire2(81, 34)    <= sub_wire176(34);
	sub_wire2(81, 35)    <= sub_wire176(35);
	sub_wire2(81, 36)    <= sub_wire176(36);
	sub_wire2(81, 37)    <= sub_wire176(37);
	sub_wire2(81, 38)    <= sub_wire176(38);
	sub_wire2(81, 39)    <= sub_wire176(39);
	sub_wire2(80, 0)    <= sub_wire177(0);
	sub_wire2(80, 1)    <= sub_wire177(1);
	sub_wire2(80, 2)    <= sub_wire177(2);
	sub_wire2(80, 3)    <= sub_wire177(3);
	sub_wire2(80, 4)    <= sub_wire177(4);
	sub_wire2(80, 5)    <= sub_wire177(5);
	sub_wire2(80, 6)    <= sub_wire177(6);
	sub_wire2(80, 7)    <= sub_wire177(7);
	sub_wire2(80, 8)    <= sub_wire177(8);
	sub_wire2(80, 9)    <= sub_wire177(9);
	sub_wire2(80, 10)    <= sub_wire177(10);
	sub_wire2(80, 11)    <= sub_wire177(11);
	sub_wire2(80, 12)    <= sub_wire177(12);
	sub_wire2(80, 13)    <= sub_wire177(13);
	sub_wire2(80, 14)    <= sub_wire177(14);
	sub_wire2(80, 15)    <= sub_wire177(15);
	sub_wire2(80, 16)    <= sub_wire177(16);
	sub_wire2(80, 17)    <= sub_wire177(17);
	sub_wire2(80, 18)    <= sub_wire177(18);
	sub_wire2(80, 19)    <= sub_wire177(19);
	sub_wire2(80, 20)    <= sub_wire177(20);
	sub_wire2(80, 21)    <= sub_wire177(21);
	sub_wire2(80, 22)    <= sub_wire177(22);
	sub_wire2(80, 23)    <= sub_wire177(23);
	sub_wire2(80, 24)    <= sub_wire177(24);
	sub_wire2(80, 25)    <= sub_wire177(25);
	sub_wire2(80, 26)    <= sub_wire177(26);
	sub_wire2(80, 27)    <= sub_wire177(27);
	sub_wire2(80, 28)    <= sub_wire177(28);
	sub_wire2(80, 29)    <= sub_wire177(29);
	sub_wire2(80, 30)    <= sub_wire177(30);
	sub_wire2(80, 31)    <= sub_wire177(31);
	sub_wire2(80, 32)    <= sub_wire177(32);
	sub_wire2(80, 33)    <= sub_wire177(33);
	sub_wire2(80, 34)    <= sub_wire177(34);
	sub_wire2(80, 35)    <= sub_wire177(35);
	sub_wire2(80, 36)    <= sub_wire177(36);
	sub_wire2(80, 37)    <= sub_wire177(37);
	sub_wire2(80, 38)    <= sub_wire177(38);
	sub_wire2(80, 39)    <= sub_wire177(39);
	sub_wire2(79, 0)    <= sub_wire178(0);
	sub_wire2(79, 1)    <= sub_wire178(1);
	sub_wire2(79, 2)    <= sub_wire178(2);
	sub_wire2(79, 3)    <= sub_wire178(3);
	sub_wire2(79, 4)    <= sub_wire178(4);
	sub_wire2(79, 5)    <= sub_wire178(5);
	sub_wire2(79, 6)    <= sub_wire178(6);
	sub_wire2(79, 7)    <= sub_wire178(7);
	sub_wire2(79, 8)    <= sub_wire178(8);
	sub_wire2(79, 9)    <= sub_wire178(9);
	sub_wire2(79, 10)    <= sub_wire178(10);
	sub_wire2(79, 11)    <= sub_wire178(11);
	sub_wire2(79, 12)    <= sub_wire178(12);
	sub_wire2(79, 13)    <= sub_wire178(13);
	sub_wire2(79, 14)    <= sub_wire178(14);
	sub_wire2(79, 15)    <= sub_wire178(15);
	sub_wire2(79, 16)    <= sub_wire178(16);
	sub_wire2(79, 17)    <= sub_wire178(17);
	sub_wire2(79, 18)    <= sub_wire178(18);
	sub_wire2(79, 19)    <= sub_wire178(19);
	sub_wire2(79, 20)    <= sub_wire178(20);
	sub_wire2(79, 21)    <= sub_wire178(21);
	sub_wire2(79, 22)    <= sub_wire178(22);
	sub_wire2(79, 23)    <= sub_wire178(23);
	sub_wire2(79, 24)    <= sub_wire178(24);
	sub_wire2(79, 25)    <= sub_wire178(25);
	sub_wire2(79, 26)    <= sub_wire178(26);
	sub_wire2(79, 27)    <= sub_wire178(27);
	sub_wire2(79, 28)    <= sub_wire178(28);
	sub_wire2(79, 29)    <= sub_wire178(29);
	sub_wire2(79, 30)    <= sub_wire178(30);
	sub_wire2(79, 31)    <= sub_wire178(31);
	sub_wire2(79, 32)    <= sub_wire178(32);
	sub_wire2(79, 33)    <= sub_wire178(33);
	sub_wire2(79, 34)    <= sub_wire178(34);
	sub_wire2(79, 35)    <= sub_wire178(35);
	sub_wire2(79, 36)    <= sub_wire178(36);
	sub_wire2(79, 37)    <= sub_wire178(37);
	sub_wire2(79, 38)    <= sub_wire178(38);
	sub_wire2(79, 39)    <= sub_wire178(39);
	sub_wire2(78, 0)    <= sub_wire179(0);
	sub_wire2(78, 1)    <= sub_wire179(1);
	sub_wire2(78, 2)    <= sub_wire179(2);
	sub_wire2(78, 3)    <= sub_wire179(3);
	sub_wire2(78, 4)    <= sub_wire179(4);
	sub_wire2(78, 5)    <= sub_wire179(5);
	sub_wire2(78, 6)    <= sub_wire179(6);
	sub_wire2(78, 7)    <= sub_wire179(7);
	sub_wire2(78, 8)    <= sub_wire179(8);
	sub_wire2(78, 9)    <= sub_wire179(9);
	sub_wire2(78, 10)    <= sub_wire179(10);
	sub_wire2(78, 11)    <= sub_wire179(11);
	sub_wire2(78, 12)    <= sub_wire179(12);
	sub_wire2(78, 13)    <= sub_wire179(13);
	sub_wire2(78, 14)    <= sub_wire179(14);
	sub_wire2(78, 15)    <= sub_wire179(15);
	sub_wire2(78, 16)    <= sub_wire179(16);
	sub_wire2(78, 17)    <= sub_wire179(17);
	sub_wire2(78, 18)    <= sub_wire179(18);
	sub_wire2(78, 19)    <= sub_wire179(19);
	sub_wire2(78, 20)    <= sub_wire179(20);
	sub_wire2(78, 21)    <= sub_wire179(21);
	sub_wire2(78, 22)    <= sub_wire179(22);
	sub_wire2(78, 23)    <= sub_wire179(23);
	sub_wire2(78, 24)    <= sub_wire179(24);
	sub_wire2(78, 25)    <= sub_wire179(25);
	sub_wire2(78, 26)    <= sub_wire179(26);
	sub_wire2(78, 27)    <= sub_wire179(27);
	sub_wire2(78, 28)    <= sub_wire179(28);
	sub_wire2(78, 29)    <= sub_wire179(29);
	sub_wire2(78, 30)    <= sub_wire179(30);
	sub_wire2(78, 31)    <= sub_wire179(31);
	sub_wire2(78, 32)    <= sub_wire179(32);
	sub_wire2(78, 33)    <= sub_wire179(33);
	sub_wire2(78, 34)    <= sub_wire179(34);
	sub_wire2(78, 35)    <= sub_wire179(35);
	sub_wire2(78, 36)    <= sub_wire179(36);
	sub_wire2(78, 37)    <= sub_wire179(37);
	sub_wire2(78, 38)    <= sub_wire179(38);
	sub_wire2(78, 39)    <= sub_wire179(39);
	sub_wire2(77, 0)    <= sub_wire180(0);
	sub_wire2(77, 1)    <= sub_wire180(1);
	sub_wire2(77, 2)    <= sub_wire180(2);
	sub_wire2(77, 3)    <= sub_wire180(3);
	sub_wire2(77, 4)    <= sub_wire180(4);
	sub_wire2(77, 5)    <= sub_wire180(5);
	sub_wire2(77, 6)    <= sub_wire180(6);
	sub_wire2(77, 7)    <= sub_wire180(7);
	sub_wire2(77, 8)    <= sub_wire180(8);
	sub_wire2(77, 9)    <= sub_wire180(9);
	sub_wire2(77, 10)    <= sub_wire180(10);
	sub_wire2(77, 11)    <= sub_wire180(11);
	sub_wire2(77, 12)    <= sub_wire180(12);
	sub_wire2(77, 13)    <= sub_wire180(13);
	sub_wire2(77, 14)    <= sub_wire180(14);
	sub_wire2(77, 15)    <= sub_wire180(15);
	sub_wire2(77, 16)    <= sub_wire180(16);
	sub_wire2(77, 17)    <= sub_wire180(17);
	sub_wire2(77, 18)    <= sub_wire180(18);
	sub_wire2(77, 19)    <= sub_wire180(19);
	sub_wire2(77, 20)    <= sub_wire180(20);
	sub_wire2(77, 21)    <= sub_wire180(21);
	sub_wire2(77, 22)    <= sub_wire180(22);
	sub_wire2(77, 23)    <= sub_wire180(23);
	sub_wire2(77, 24)    <= sub_wire180(24);
	sub_wire2(77, 25)    <= sub_wire180(25);
	sub_wire2(77, 26)    <= sub_wire180(26);
	sub_wire2(77, 27)    <= sub_wire180(27);
	sub_wire2(77, 28)    <= sub_wire180(28);
	sub_wire2(77, 29)    <= sub_wire180(29);
	sub_wire2(77, 30)    <= sub_wire180(30);
	sub_wire2(77, 31)    <= sub_wire180(31);
	sub_wire2(77, 32)    <= sub_wire180(32);
	sub_wire2(77, 33)    <= sub_wire180(33);
	sub_wire2(77, 34)    <= sub_wire180(34);
	sub_wire2(77, 35)    <= sub_wire180(35);
	sub_wire2(77, 36)    <= sub_wire180(36);
	sub_wire2(77, 37)    <= sub_wire180(37);
	sub_wire2(77, 38)    <= sub_wire180(38);
	sub_wire2(77, 39)    <= sub_wire180(39);
	sub_wire2(76, 0)    <= sub_wire181(0);
	sub_wire2(76, 1)    <= sub_wire181(1);
	sub_wire2(76, 2)    <= sub_wire181(2);
	sub_wire2(76, 3)    <= sub_wire181(3);
	sub_wire2(76, 4)    <= sub_wire181(4);
	sub_wire2(76, 5)    <= sub_wire181(5);
	sub_wire2(76, 6)    <= sub_wire181(6);
	sub_wire2(76, 7)    <= sub_wire181(7);
	sub_wire2(76, 8)    <= sub_wire181(8);
	sub_wire2(76, 9)    <= sub_wire181(9);
	sub_wire2(76, 10)    <= sub_wire181(10);
	sub_wire2(76, 11)    <= sub_wire181(11);
	sub_wire2(76, 12)    <= sub_wire181(12);
	sub_wire2(76, 13)    <= sub_wire181(13);
	sub_wire2(76, 14)    <= sub_wire181(14);
	sub_wire2(76, 15)    <= sub_wire181(15);
	sub_wire2(76, 16)    <= sub_wire181(16);
	sub_wire2(76, 17)    <= sub_wire181(17);
	sub_wire2(76, 18)    <= sub_wire181(18);
	sub_wire2(76, 19)    <= sub_wire181(19);
	sub_wire2(76, 20)    <= sub_wire181(20);
	sub_wire2(76, 21)    <= sub_wire181(21);
	sub_wire2(76, 22)    <= sub_wire181(22);
	sub_wire2(76, 23)    <= sub_wire181(23);
	sub_wire2(76, 24)    <= sub_wire181(24);
	sub_wire2(76, 25)    <= sub_wire181(25);
	sub_wire2(76, 26)    <= sub_wire181(26);
	sub_wire2(76, 27)    <= sub_wire181(27);
	sub_wire2(76, 28)    <= sub_wire181(28);
	sub_wire2(76, 29)    <= sub_wire181(29);
	sub_wire2(76, 30)    <= sub_wire181(30);
	sub_wire2(76, 31)    <= sub_wire181(31);
	sub_wire2(76, 32)    <= sub_wire181(32);
	sub_wire2(76, 33)    <= sub_wire181(33);
	sub_wire2(76, 34)    <= sub_wire181(34);
	sub_wire2(76, 35)    <= sub_wire181(35);
	sub_wire2(76, 36)    <= sub_wire181(36);
	sub_wire2(76, 37)    <= sub_wire181(37);
	sub_wire2(76, 38)    <= sub_wire181(38);
	sub_wire2(76, 39)    <= sub_wire181(39);
	sub_wire2(75, 0)    <= sub_wire182(0);
	sub_wire2(75, 1)    <= sub_wire182(1);
	sub_wire2(75, 2)    <= sub_wire182(2);
	sub_wire2(75, 3)    <= sub_wire182(3);
	sub_wire2(75, 4)    <= sub_wire182(4);
	sub_wire2(75, 5)    <= sub_wire182(5);
	sub_wire2(75, 6)    <= sub_wire182(6);
	sub_wire2(75, 7)    <= sub_wire182(7);
	sub_wire2(75, 8)    <= sub_wire182(8);
	sub_wire2(75, 9)    <= sub_wire182(9);
	sub_wire2(75, 10)    <= sub_wire182(10);
	sub_wire2(75, 11)    <= sub_wire182(11);
	sub_wire2(75, 12)    <= sub_wire182(12);
	sub_wire2(75, 13)    <= sub_wire182(13);
	sub_wire2(75, 14)    <= sub_wire182(14);
	sub_wire2(75, 15)    <= sub_wire182(15);
	sub_wire2(75, 16)    <= sub_wire182(16);
	sub_wire2(75, 17)    <= sub_wire182(17);
	sub_wire2(75, 18)    <= sub_wire182(18);
	sub_wire2(75, 19)    <= sub_wire182(19);
	sub_wire2(75, 20)    <= sub_wire182(20);
	sub_wire2(75, 21)    <= sub_wire182(21);
	sub_wire2(75, 22)    <= sub_wire182(22);
	sub_wire2(75, 23)    <= sub_wire182(23);
	sub_wire2(75, 24)    <= sub_wire182(24);
	sub_wire2(75, 25)    <= sub_wire182(25);
	sub_wire2(75, 26)    <= sub_wire182(26);
	sub_wire2(75, 27)    <= sub_wire182(27);
	sub_wire2(75, 28)    <= sub_wire182(28);
	sub_wire2(75, 29)    <= sub_wire182(29);
	sub_wire2(75, 30)    <= sub_wire182(30);
	sub_wire2(75, 31)    <= sub_wire182(31);
	sub_wire2(75, 32)    <= sub_wire182(32);
	sub_wire2(75, 33)    <= sub_wire182(33);
	sub_wire2(75, 34)    <= sub_wire182(34);
	sub_wire2(75, 35)    <= sub_wire182(35);
	sub_wire2(75, 36)    <= sub_wire182(36);
	sub_wire2(75, 37)    <= sub_wire182(37);
	sub_wire2(75, 38)    <= sub_wire182(38);
	sub_wire2(75, 39)    <= sub_wire182(39);
	sub_wire2(74, 0)    <= sub_wire183(0);
	sub_wire2(74, 1)    <= sub_wire183(1);
	sub_wire2(74, 2)    <= sub_wire183(2);
	sub_wire2(74, 3)    <= sub_wire183(3);
	sub_wire2(74, 4)    <= sub_wire183(4);
	sub_wire2(74, 5)    <= sub_wire183(5);
	sub_wire2(74, 6)    <= sub_wire183(6);
	sub_wire2(74, 7)    <= sub_wire183(7);
	sub_wire2(74, 8)    <= sub_wire183(8);
	sub_wire2(74, 9)    <= sub_wire183(9);
	sub_wire2(74, 10)    <= sub_wire183(10);
	sub_wire2(74, 11)    <= sub_wire183(11);
	sub_wire2(74, 12)    <= sub_wire183(12);
	sub_wire2(74, 13)    <= sub_wire183(13);
	sub_wire2(74, 14)    <= sub_wire183(14);
	sub_wire2(74, 15)    <= sub_wire183(15);
	sub_wire2(74, 16)    <= sub_wire183(16);
	sub_wire2(74, 17)    <= sub_wire183(17);
	sub_wire2(74, 18)    <= sub_wire183(18);
	sub_wire2(74, 19)    <= sub_wire183(19);
	sub_wire2(74, 20)    <= sub_wire183(20);
	sub_wire2(74, 21)    <= sub_wire183(21);
	sub_wire2(74, 22)    <= sub_wire183(22);
	sub_wire2(74, 23)    <= sub_wire183(23);
	sub_wire2(74, 24)    <= sub_wire183(24);
	sub_wire2(74, 25)    <= sub_wire183(25);
	sub_wire2(74, 26)    <= sub_wire183(26);
	sub_wire2(74, 27)    <= sub_wire183(27);
	sub_wire2(74, 28)    <= sub_wire183(28);
	sub_wire2(74, 29)    <= sub_wire183(29);
	sub_wire2(74, 30)    <= sub_wire183(30);
	sub_wire2(74, 31)    <= sub_wire183(31);
	sub_wire2(74, 32)    <= sub_wire183(32);
	sub_wire2(74, 33)    <= sub_wire183(33);
	sub_wire2(74, 34)    <= sub_wire183(34);
	sub_wire2(74, 35)    <= sub_wire183(35);
	sub_wire2(74, 36)    <= sub_wire183(36);
	sub_wire2(74, 37)    <= sub_wire183(37);
	sub_wire2(74, 38)    <= sub_wire183(38);
	sub_wire2(74, 39)    <= sub_wire183(39);
	sub_wire2(73, 0)    <= sub_wire184(0);
	sub_wire2(73, 1)    <= sub_wire184(1);
	sub_wire2(73, 2)    <= sub_wire184(2);
	sub_wire2(73, 3)    <= sub_wire184(3);
	sub_wire2(73, 4)    <= sub_wire184(4);
	sub_wire2(73, 5)    <= sub_wire184(5);
	sub_wire2(73, 6)    <= sub_wire184(6);
	sub_wire2(73, 7)    <= sub_wire184(7);
	sub_wire2(73, 8)    <= sub_wire184(8);
	sub_wire2(73, 9)    <= sub_wire184(9);
	sub_wire2(73, 10)    <= sub_wire184(10);
	sub_wire2(73, 11)    <= sub_wire184(11);
	sub_wire2(73, 12)    <= sub_wire184(12);
	sub_wire2(73, 13)    <= sub_wire184(13);
	sub_wire2(73, 14)    <= sub_wire184(14);
	sub_wire2(73, 15)    <= sub_wire184(15);
	sub_wire2(73, 16)    <= sub_wire184(16);
	sub_wire2(73, 17)    <= sub_wire184(17);
	sub_wire2(73, 18)    <= sub_wire184(18);
	sub_wire2(73, 19)    <= sub_wire184(19);
	sub_wire2(73, 20)    <= sub_wire184(20);
	sub_wire2(73, 21)    <= sub_wire184(21);
	sub_wire2(73, 22)    <= sub_wire184(22);
	sub_wire2(73, 23)    <= sub_wire184(23);
	sub_wire2(73, 24)    <= sub_wire184(24);
	sub_wire2(73, 25)    <= sub_wire184(25);
	sub_wire2(73, 26)    <= sub_wire184(26);
	sub_wire2(73, 27)    <= sub_wire184(27);
	sub_wire2(73, 28)    <= sub_wire184(28);
	sub_wire2(73, 29)    <= sub_wire184(29);
	sub_wire2(73, 30)    <= sub_wire184(30);
	sub_wire2(73, 31)    <= sub_wire184(31);
	sub_wire2(73, 32)    <= sub_wire184(32);
	sub_wire2(73, 33)    <= sub_wire184(33);
	sub_wire2(73, 34)    <= sub_wire184(34);
	sub_wire2(73, 35)    <= sub_wire184(35);
	sub_wire2(73, 36)    <= sub_wire184(36);
	sub_wire2(73, 37)    <= sub_wire184(37);
	sub_wire2(73, 38)    <= sub_wire184(38);
	sub_wire2(73, 39)    <= sub_wire184(39);
	sub_wire2(72, 0)    <= sub_wire185(0);
	sub_wire2(72, 1)    <= sub_wire185(1);
	sub_wire2(72, 2)    <= sub_wire185(2);
	sub_wire2(72, 3)    <= sub_wire185(3);
	sub_wire2(72, 4)    <= sub_wire185(4);
	sub_wire2(72, 5)    <= sub_wire185(5);
	sub_wire2(72, 6)    <= sub_wire185(6);
	sub_wire2(72, 7)    <= sub_wire185(7);
	sub_wire2(72, 8)    <= sub_wire185(8);
	sub_wire2(72, 9)    <= sub_wire185(9);
	sub_wire2(72, 10)    <= sub_wire185(10);
	sub_wire2(72, 11)    <= sub_wire185(11);
	sub_wire2(72, 12)    <= sub_wire185(12);
	sub_wire2(72, 13)    <= sub_wire185(13);
	sub_wire2(72, 14)    <= sub_wire185(14);
	sub_wire2(72, 15)    <= sub_wire185(15);
	sub_wire2(72, 16)    <= sub_wire185(16);
	sub_wire2(72, 17)    <= sub_wire185(17);
	sub_wire2(72, 18)    <= sub_wire185(18);
	sub_wire2(72, 19)    <= sub_wire185(19);
	sub_wire2(72, 20)    <= sub_wire185(20);
	sub_wire2(72, 21)    <= sub_wire185(21);
	sub_wire2(72, 22)    <= sub_wire185(22);
	sub_wire2(72, 23)    <= sub_wire185(23);
	sub_wire2(72, 24)    <= sub_wire185(24);
	sub_wire2(72, 25)    <= sub_wire185(25);
	sub_wire2(72, 26)    <= sub_wire185(26);
	sub_wire2(72, 27)    <= sub_wire185(27);
	sub_wire2(72, 28)    <= sub_wire185(28);
	sub_wire2(72, 29)    <= sub_wire185(29);
	sub_wire2(72, 30)    <= sub_wire185(30);
	sub_wire2(72, 31)    <= sub_wire185(31);
	sub_wire2(72, 32)    <= sub_wire185(32);
	sub_wire2(72, 33)    <= sub_wire185(33);
	sub_wire2(72, 34)    <= sub_wire185(34);
	sub_wire2(72, 35)    <= sub_wire185(35);
	sub_wire2(72, 36)    <= sub_wire185(36);
	sub_wire2(72, 37)    <= sub_wire185(37);
	sub_wire2(72, 38)    <= sub_wire185(38);
	sub_wire2(72, 39)    <= sub_wire185(39);
	sub_wire2(71, 0)    <= sub_wire186(0);
	sub_wire2(71, 1)    <= sub_wire186(1);
	sub_wire2(71, 2)    <= sub_wire186(2);
	sub_wire2(71, 3)    <= sub_wire186(3);
	sub_wire2(71, 4)    <= sub_wire186(4);
	sub_wire2(71, 5)    <= sub_wire186(5);
	sub_wire2(71, 6)    <= sub_wire186(6);
	sub_wire2(71, 7)    <= sub_wire186(7);
	sub_wire2(71, 8)    <= sub_wire186(8);
	sub_wire2(71, 9)    <= sub_wire186(9);
	sub_wire2(71, 10)    <= sub_wire186(10);
	sub_wire2(71, 11)    <= sub_wire186(11);
	sub_wire2(71, 12)    <= sub_wire186(12);
	sub_wire2(71, 13)    <= sub_wire186(13);
	sub_wire2(71, 14)    <= sub_wire186(14);
	sub_wire2(71, 15)    <= sub_wire186(15);
	sub_wire2(71, 16)    <= sub_wire186(16);
	sub_wire2(71, 17)    <= sub_wire186(17);
	sub_wire2(71, 18)    <= sub_wire186(18);
	sub_wire2(71, 19)    <= sub_wire186(19);
	sub_wire2(71, 20)    <= sub_wire186(20);
	sub_wire2(71, 21)    <= sub_wire186(21);
	sub_wire2(71, 22)    <= sub_wire186(22);
	sub_wire2(71, 23)    <= sub_wire186(23);
	sub_wire2(71, 24)    <= sub_wire186(24);
	sub_wire2(71, 25)    <= sub_wire186(25);
	sub_wire2(71, 26)    <= sub_wire186(26);
	sub_wire2(71, 27)    <= sub_wire186(27);
	sub_wire2(71, 28)    <= sub_wire186(28);
	sub_wire2(71, 29)    <= sub_wire186(29);
	sub_wire2(71, 30)    <= sub_wire186(30);
	sub_wire2(71, 31)    <= sub_wire186(31);
	sub_wire2(71, 32)    <= sub_wire186(32);
	sub_wire2(71, 33)    <= sub_wire186(33);
	sub_wire2(71, 34)    <= sub_wire186(34);
	sub_wire2(71, 35)    <= sub_wire186(35);
	sub_wire2(71, 36)    <= sub_wire186(36);
	sub_wire2(71, 37)    <= sub_wire186(37);
	sub_wire2(71, 38)    <= sub_wire186(38);
	sub_wire2(71, 39)    <= sub_wire186(39);
	sub_wire2(70, 0)    <= sub_wire187(0);
	sub_wire2(70, 1)    <= sub_wire187(1);
	sub_wire2(70, 2)    <= sub_wire187(2);
	sub_wire2(70, 3)    <= sub_wire187(3);
	sub_wire2(70, 4)    <= sub_wire187(4);
	sub_wire2(70, 5)    <= sub_wire187(5);
	sub_wire2(70, 6)    <= sub_wire187(6);
	sub_wire2(70, 7)    <= sub_wire187(7);
	sub_wire2(70, 8)    <= sub_wire187(8);
	sub_wire2(70, 9)    <= sub_wire187(9);
	sub_wire2(70, 10)    <= sub_wire187(10);
	sub_wire2(70, 11)    <= sub_wire187(11);
	sub_wire2(70, 12)    <= sub_wire187(12);
	sub_wire2(70, 13)    <= sub_wire187(13);
	sub_wire2(70, 14)    <= sub_wire187(14);
	sub_wire2(70, 15)    <= sub_wire187(15);
	sub_wire2(70, 16)    <= sub_wire187(16);
	sub_wire2(70, 17)    <= sub_wire187(17);
	sub_wire2(70, 18)    <= sub_wire187(18);
	sub_wire2(70, 19)    <= sub_wire187(19);
	sub_wire2(70, 20)    <= sub_wire187(20);
	sub_wire2(70, 21)    <= sub_wire187(21);
	sub_wire2(70, 22)    <= sub_wire187(22);
	sub_wire2(70, 23)    <= sub_wire187(23);
	sub_wire2(70, 24)    <= sub_wire187(24);
	sub_wire2(70, 25)    <= sub_wire187(25);
	sub_wire2(70, 26)    <= sub_wire187(26);
	sub_wire2(70, 27)    <= sub_wire187(27);
	sub_wire2(70, 28)    <= sub_wire187(28);
	sub_wire2(70, 29)    <= sub_wire187(29);
	sub_wire2(70, 30)    <= sub_wire187(30);
	sub_wire2(70, 31)    <= sub_wire187(31);
	sub_wire2(70, 32)    <= sub_wire187(32);
	sub_wire2(70, 33)    <= sub_wire187(33);
	sub_wire2(70, 34)    <= sub_wire187(34);
	sub_wire2(70, 35)    <= sub_wire187(35);
	sub_wire2(70, 36)    <= sub_wire187(36);
	sub_wire2(70, 37)    <= sub_wire187(37);
	sub_wire2(70, 38)    <= sub_wire187(38);
	sub_wire2(70, 39)    <= sub_wire187(39);
	sub_wire2(69, 0)    <= sub_wire188(0);
	sub_wire2(69, 1)    <= sub_wire188(1);
	sub_wire2(69, 2)    <= sub_wire188(2);
	sub_wire2(69, 3)    <= sub_wire188(3);
	sub_wire2(69, 4)    <= sub_wire188(4);
	sub_wire2(69, 5)    <= sub_wire188(5);
	sub_wire2(69, 6)    <= sub_wire188(6);
	sub_wire2(69, 7)    <= sub_wire188(7);
	sub_wire2(69, 8)    <= sub_wire188(8);
	sub_wire2(69, 9)    <= sub_wire188(9);
	sub_wire2(69, 10)    <= sub_wire188(10);
	sub_wire2(69, 11)    <= sub_wire188(11);
	sub_wire2(69, 12)    <= sub_wire188(12);
	sub_wire2(69, 13)    <= sub_wire188(13);
	sub_wire2(69, 14)    <= sub_wire188(14);
	sub_wire2(69, 15)    <= sub_wire188(15);
	sub_wire2(69, 16)    <= sub_wire188(16);
	sub_wire2(69, 17)    <= sub_wire188(17);
	sub_wire2(69, 18)    <= sub_wire188(18);
	sub_wire2(69, 19)    <= sub_wire188(19);
	sub_wire2(69, 20)    <= sub_wire188(20);
	sub_wire2(69, 21)    <= sub_wire188(21);
	sub_wire2(69, 22)    <= sub_wire188(22);
	sub_wire2(69, 23)    <= sub_wire188(23);
	sub_wire2(69, 24)    <= sub_wire188(24);
	sub_wire2(69, 25)    <= sub_wire188(25);
	sub_wire2(69, 26)    <= sub_wire188(26);
	sub_wire2(69, 27)    <= sub_wire188(27);
	sub_wire2(69, 28)    <= sub_wire188(28);
	sub_wire2(69, 29)    <= sub_wire188(29);
	sub_wire2(69, 30)    <= sub_wire188(30);
	sub_wire2(69, 31)    <= sub_wire188(31);
	sub_wire2(69, 32)    <= sub_wire188(32);
	sub_wire2(69, 33)    <= sub_wire188(33);
	sub_wire2(69, 34)    <= sub_wire188(34);
	sub_wire2(69, 35)    <= sub_wire188(35);
	sub_wire2(69, 36)    <= sub_wire188(36);
	sub_wire2(69, 37)    <= sub_wire188(37);
	sub_wire2(69, 38)    <= sub_wire188(38);
	sub_wire2(69, 39)    <= sub_wire188(39);
	sub_wire2(68, 0)    <= sub_wire189(0);
	sub_wire2(68, 1)    <= sub_wire189(1);
	sub_wire2(68, 2)    <= sub_wire189(2);
	sub_wire2(68, 3)    <= sub_wire189(3);
	sub_wire2(68, 4)    <= sub_wire189(4);
	sub_wire2(68, 5)    <= sub_wire189(5);
	sub_wire2(68, 6)    <= sub_wire189(6);
	sub_wire2(68, 7)    <= sub_wire189(7);
	sub_wire2(68, 8)    <= sub_wire189(8);
	sub_wire2(68, 9)    <= sub_wire189(9);
	sub_wire2(68, 10)    <= sub_wire189(10);
	sub_wire2(68, 11)    <= sub_wire189(11);
	sub_wire2(68, 12)    <= sub_wire189(12);
	sub_wire2(68, 13)    <= sub_wire189(13);
	sub_wire2(68, 14)    <= sub_wire189(14);
	sub_wire2(68, 15)    <= sub_wire189(15);
	sub_wire2(68, 16)    <= sub_wire189(16);
	sub_wire2(68, 17)    <= sub_wire189(17);
	sub_wire2(68, 18)    <= sub_wire189(18);
	sub_wire2(68, 19)    <= sub_wire189(19);
	sub_wire2(68, 20)    <= sub_wire189(20);
	sub_wire2(68, 21)    <= sub_wire189(21);
	sub_wire2(68, 22)    <= sub_wire189(22);
	sub_wire2(68, 23)    <= sub_wire189(23);
	sub_wire2(68, 24)    <= sub_wire189(24);
	sub_wire2(68, 25)    <= sub_wire189(25);
	sub_wire2(68, 26)    <= sub_wire189(26);
	sub_wire2(68, 27)    <= sub_wire189(27);
	sub_wire2(68, 28)    <= sub_wire189(28);
	sub_wire2(68, 29)    <= sub_wire189(29);
	sub_wire2(68, 30)    <= sub_wire189(30);
	sub_wire2(68, 31)    <= sub_wire189(31);
	sub_wire2(68, 32)    <= sub_wire189(32);
	sub_wire2(68, 33)    <= sub_wire189(33);
	sub_wire2(68, 34)    <= sub_wire189(34);
	sub_wire2(68, 35)    <= sub_wire189(35);
	sub_wire2(68, 36)    <= sub_wire189(36);
	sub_wire2(68, 37)    <= sub_wire189(37);
	sub_wire2(68, 38)    <= sub_wire189(38);
	sub_wire2(68, 39)    <= sub_wire189(39);
	sub_wire2(67, 0)    <= sub_wire190(0);
	sub_wire2(67, 1)    <= sub_wire190(1);
	sub_wire2(67, 2)    <= sub_wire190(2);
	sub_wire2(67, 3)    <= sub_wire190(3);
	sub_wire2(67, 4)    <= sub_wire190(4);
	sub_wire2(67, 5)    <= sub_wire190(5);
	sub_wire2(67, 6)    <= sub_wire190(6);
	sub_wire2(67, 7)    <= sub_wire190(7);
	sub_wire2(67, 8)    <= sub_wire190(8);
	sub_wire2(67, 9)    <= sub_wire190(9);
	sub_wire2(67, 10)    <= sub_wire190(10);
	sub_wire2(67, 11)    <= sub_wire190(11);
	sub_wire2(67, 12)    <= sub_wire190(12);
	sub_wire2(67, 13)    <= sub_wire190(13);
	sub_wire2(67, 14)    <= sub_wire190(14);
	sub_wire2(67, 15)    <= sub_wire190(15);
	sub_wire2(67, 16)    <= sub_wire190(16);
	sub_wire2(67, 17)    <= sub_wire190(17);
	sub_wire2(67, 18)    <= sub_wire190(18);
	sub_wire2(67, 19)    <= sub_wire190(19);
	sub_wire2(67, 20)    <= sub_wire190(20);
	sub_wire2(67, 21)    <= sub_wire190(21);
	sub_wire2(67, 22)    <= sub_wire190(22);
	sub_wire2(67, 23)    <= sub_wire190(23);
	sub_wire2(67, 24)    <= sub_wire190(24);
	sub_wire2(67, 25)    <= sub_wire190(25);
	sub_wire2(67, 26)    <= sub_wire190(26);
	sub_wire2(67, 27)    <= sub_wire190(27);
	sub_wire2(67, 28)    <= sub_wire190(28);
	sub_wire2(67, 29)    <= sub_wire190(29);
	sub_wire2(67, 30)    <= sub_wire190(30);
	sub_wire2(67, 31)    <= sub_wire190(31);
	sub_wire2(67, 32)    <= sub_wire190(32);
	sub_wire2(67, 33)    <= sub_wire190(33);
	sub_wire2(67, 34)    <= sub_wire190(34);
	sub_wire2(67, 35)    <= sub_wire190(35);
	sub_wire2(67, 36)    <= sub_wire190(36);
	sub_wire2(67, 37)    <= sub_wire190(37);
	sub_wire2(67, 38)    <= sub_wire190(38);
	sub_wire2(67, 39)    <= sub_wire190(39);
	sub_wire2(66, 0)    <= sub_wire191(0);
	sub_wire2(66, 1)    <= sub_wire191(1);
	sub_wire2(66, 2)    <= sub_wire191(2);
	sub_wire2(66, 3)    <= sub_wire191(3);
	sub_wire2(66, 4)    <= sub_wire191(4);
	sub_wire2(66, 5)    <= sub_wire191(5);
	sub_wire2(66, 6)    <= sub_wire191(6);
	sub_wire2(66, 7)    <= sub_wire191(7);
	sub_wire2(66, 8)    <= sub_wire191(8);
	sub_wire2(66, 9)    <= sub_wire191(9);
	sub_wire2(66, 10)    <= sub_wire191(10);
	sub_wire2(66, 11)    <= sub_wire191(11);
	sub_wire2(66, 12)    <= sub_wire191(12);
	sub_wire2(66, 13)    <= sub_wire191(13);
	sub_wire2(66, 14)    <= sub_wire191(14);
	sub_wire2(66, 15)    <= sub_wire191(15);
	sub_wire2(66, 16)    <= sub_wire191(16);
	sub_wire2(66, 17)    <= sub_wire191(17);
	sub_wire2(66, 18)    <= sub_wire191(18);
	sub_wire2(66, 19)    <= sub_wire191(19);
	sub_wire2(66, 20)    <= sub_wire191(20);
	sub_wire2(66, 21)    <= sub_wire191(21);
	sub_wire2(66, 22)    <= sub_wire191(22);
	sub_wire2(66, 23)    <= sub_wire191(23);
	sub_wire2(66, 24)    <= sub_wire191(24);
	sub_wire2(66, 25)    <= sub_wire191(25);
	sub_wire2(66, 26)    <= sub_wire191(26);
	sub_wire2(66, 27)    <= sub_wire191(27);
	sub_wire2(66, 28)    <= sub_wire191(28);
	sub_wire2(66, 29)    <= sub_wire191(29);
	sub_wire2(66, 30)    <= sub_wire191(30);
	sub_wire2(66, 31)    <= sub_wire191(31);
	sub_wire2(66, 32)    <= sub_wire191(32);
	sub_wire2(66, 33)    <= sub_wire191(33);
	sub_wire2(66, 34)    <= sub_wire191(34);
	sub_wire2(66, 35)    <= sub_wire191(35);
	sub_wire2(66, 36)    <= sub_wire191(36);
	sub_wire2(66, 37)    <= sub_wire191(37);
	sub_wire2(66, 38)    <= sub_wire191(38);
	sub_wire2(66, 39)    <= sub_wire191(39);
	sub_wire2(65, 0)    <= sub_wire192(0);
	sub_wire2(65, 1)    <= sub_wire192(1);
	sub_wire2(65, 2)    <= sub_wire192(2);
	sub_wire2(65, 3)    <= sub_wire192(3);
	sub_wire2(65, 4)    <= sub_wire192(4);
	sub_wire2(65, 5)    <= sub_wire192(5);
	sub_wire2(65, 6)    <= sub_wire192(6);
	sub_wire2(65, 7)    <= sub_wire192(7);
	sub_wire2(65, 8)    <= sub_wire192(8);
	sub_wire2(65, 9)    <= sub_wire192(9);
	sub_wire2(65, 10)    <= sub_wire192(10);
	sub_wire2(65, 11)    <= sub_wire192(11);
	sub_wire2(65, 12)    <= sub_wire192(12);
	sub_wire2(65, 13)    <= sub_wire192(13);
	sub_wire2(65, 14)    <= sub_wire192(14);
	sub_wire2(65, 15)    <= sub_wire192(15);
	sub_wire2(65, 16)    <= sub_wire192(16);
	sub_wire2(65, 17)    <= sub_wire192(17);
	sub_wire2(65, 18)    <= sub_wire192(18);
	sub_wire2(65, 19)    <= sub_wire192(19);
	sub_wire2(65, 20)    <= sub_wire192(20);
	sub_wire2(65, 21)    <= sub_wire192(21);
	sub_wire2(65, 22)    <= sub_wire192(22);
	sub_wire2(65, 23)    <= sub_wire192(23);
	sub_wire2(65, 24)    <= sub_wire192(24);
	sub_wire2(65, 25)    <= sub_wire192(25);
	sub_wire2(65, 26)    <= sub_wire192(26);
	sub_wire2(65, 27)    <= sub_wire192(27);
	sub_wire2(65, 28)    <= sub_wire192(28);
	sub_wire2(65, 29)    <= sub_wire192(29);
	sub_wire2(65, 30)    <= sub_wire192(30);
	sub_wire2(65, 31)    <= sub_wire192(31);
	sub_wire2(65, 32)    <= sub_wire192(32);
	sub_wire2(65, 33)    <= sub_wire192(33);
	sub_wire2(65, 34)    <= sub_wire192(34);
	sub_wire2(65, 35)    <= sub_wire192(35);
	sub_wire2(65, 36)    <= sub_wire192(36);
	sub_wire2(65, 37)    <= sub_wire192(37);
	sub_wire2(65, 38)    <= sub_wire192(38);
	sub_wire2(65, 39)    <= sub_wire192(39);
	sub_wire2(64, 0)    <= sub_wire193(0);
	sub_wire2(64, 1)    <= sub_wire193(1);
	sub_wire2(64, 2)    <= sub_wire193(2);
	sub_wire2(64, 3)    <= sub_wire193(3);
	sub_wire2(64, 4)    <= sub_wire193(4);
	sub_wire2(64, 5)    <= sub_wire193(5);
	sub_wire2(64, 6)    <= sub_wire193(6);
	sub_wire2(64, 7)    <= sub_wire193(7);
	sub_wire2(64, 8)    <= sub_wire193(8);
	sub_wire2(64, 9)    <= sub_wire193(9);
	sub_wire2(64, 10)    <= sub_wire193(10);
	sub_wire2(64, 11)    <= sub_wire193(11);
	sub_wire2(64, 12)    <= sub_wire193(12);
	sub_wire2(64, 13)    <= sub_wire193(13);
	sub_wire2(64, 14)    <= sub_wire193(14);
	sub_wire2(64, 15)    <= sub_wire193(15);
	sub_wire2(64, 16)    <= sub_wire193(16);
	sub_wire2(64, 17)    <= sub_wire193(17);
	sub_wire2(64, 18)    <= sub_wire193(18);
	sub_wire2(64, 19)    <= sub_wire193(19);
	sub_wire2(64, 20)    <= sub_wire193(20);
	sub_wire2(64, 21)    <= sub_wire193(21);
	sub_wire2(64, 22)    <= sub_wire193(22);
	sub_wire2(64, 23)    <= sub_wire193(23);
	sub_wire2(64, 24)    <= sub_wire193(24);
	sub_wire2(64, 25)    <= sub_wire193(25);
	sub_wire2(64, 26)    <= sub_wire193(26);
	sub_wire2(64, 27)    <= sub_wire193(27);
	sub_wire2(64, 28)    <= sub_wire193(28);
	sub_wire2(64, 29)    <= sub_wire193(29);
	sub_wire2(64, 30)    <= sub_wire193(30);
	sub_wire2(64, 31)    <= sub_wire193(31);
	sub_wire2(64, 32)    <= sub_wire193(32);
	sub_wire2(64, 33)    <= sub_wire193(33);
	sub_wire2(64, 34)    <= sub_wire193(34);
	sub_wire2(64, 35)    <= sub_wire193(35);
	sub_wire2(64, 36)    <= sub_wire193(36);
	sub_wire2(64, 37)    <= sub_wire193(37);
	sub_wire2(64, 38)    <= sub_wire193(38);
	sub_wire2(64, 39)    <= sub_wire193(39);
	sub_wire2(63, 0)    <= sub_wire194(0);
	sub_wire2(63, 1)    <= sub_wire194(1);
	sub_wire2(63, 2)    <= sub_wire194(2);
	sub_wire2(63, 3)    <= sub_wire194(3);
	sub_wire2(63, 4)    <= sub_wire194(4);
	sub_wire2(63, 5)    <= sub_wire194(5);
	sub_wire2(63, 6)    <= sub_wire194(6);
	sub_wire2(63, 7)    <= sub_wire194(7);
	sub_wire2(63, 8)    <= sub_wire194(8);
	sub_wire2(63, 9)    <= sub_wire194(9);
	sub_wire2(63, 10)    <= sub_wire194(10);
	sub_wire2(63, 11)    <= sub_wire194(11);
	sub_wire2(63, 12)    <= sub_wire194(12);
	sub_wire2(63, 13)    <= sub_wire194(13);
	sub_wire2(63, 14)    <= sub_wire194(14);
	sub_wire2(63, 15)    <= sub_wire194(15);
	sub_wire2(63, 16)    <= sub_wire194(16);
	sub_wire2(63, 17)    <= sub_wire194(17);
	sub_wire2(63, 18)    <= sub_wire194(18);
	sub_wire2(63, 19)    <= sub_wire194(19);
	sub_wire2(63, 20)    <= sub_wire194(20);
	sub_wire2(63, 21)    <= sub_wire194(21);
	sub_wire2(63, 22)    <= sub_wire194(22);
	sub_wire2(63, 23)    <= sub_wire194(23);
	sub_wire2(63, 24)    <= sub_wire194(24);
	sub_wire2(63, 25)    <= sub_wire194(25);
	sub_wire2(63, 26)    <= sub_wire194(26);
	sub_wire2(63, 27)    <= sub_wire194(27);
	sub_wire2(63, 28)    <= sub_wire194(28);
	sub_wire2(63, 29)    <= sub_wire194(29);
	sub_wire2(63, 30)    <= sub_wire194(30);
	sub_wire2(63, 31)    <= sub_wire194(31);
	sub_wire2(63, 32)    <= sub_wire194(32);
	sub_wire2(63, 33)    <= sub_wire194(33);
	sub_wire2(63, 34)    <= sub_wire194(34);
	sub_wire2(63, 35)    <= sub_wire194(35);
	sub_wire2(63, 36)    <= sub_wire194(36);
	sub_wire2(63, 37)    <= sub_wire194(37);
	sub_wire2(63, 38)    <= sub_wire194(38);
	sub_wire2(63, 39)    <= sub_wire194(39);
	sub_wire2(62, 0)    <= sub_wire195(0);
	sub_wire2(62, 1)    <= sub_wire195(1);
	sub_wire2(62, 2)    <= sub_wire195(2);
	sub_wire2(62, 3)    <= sub_wire195(3);
	sub_wire2(62, 4)    <= sub_wire195(4);
	sub_wire2(62, 5)    <= sub_wire195(5);
	sub_wire2(62, 6)    <= sub_wire195(6);
	sub_wire2(62, 7)    <= sub_wire195(7);
	sub_wire2(62, 8)    <= sub_wire195(8);
	sub_wire2(62, 9)    <= sub_wire195(9);
	sub_wire2(62, 10)    <= sub_wire195(10);
	sub_wire2(62, 11)    <= sub_wire195(11);
	sub_wire2(62, 12)    <= sub_wire195(12);
	sub_wire2(62, 13)    <= sub_wire195(13);
	sub_wire2(62, 14)    <= sub_wire195(14);
	sub_wire2(62, 15)    <= sub_wire195(15);
	sub_wire2(62, 16)    <= sub_wire195(16);
	sub_wire2(62, 17)    <= sub_wire195(17);
	sub_wire2(62, 18)    <= sub_wire195(18);
	sub_wire2(62, 19)    <= sub_wire195(19);
	sub_wire2(62, 20)    <= sub_wire195(20);
	sub_wire2(62, 21)    <= sub_wire195(21);
	sub_wire2(62, 22)    <= sub_wire195(22);
	sub_wire2(62, 23)    <= sub_wire195(23);
	sub_wire2(62, 24)    <= sub_wire195(24);
	sub_wire2(62, 25)    <= sub_wire195(25);
	sub_wire2(62, 26)    <= sub_wire195(26);
	sub_wire2(62, 27)    <= sub_wire195(27);
	sub_wire2(62, 28)    <= sub_wire195(28);
	sub_wire2(62, 29)    <= sub_wire195(29);
	sub_wire2(62, 30)    <= sub_wire195(30);
	sub_wire2(62, 31)    <= sub_wire195(31);
	sub_wire2(62, 32)    <= sub_wire195(32);
	sub_wire2(62, 33)    <= sub_wire195(33);
	sub_wire2(62, 34)    <= sub_wire195(34);
	sub_wire2(62, 35)    <= sub_wire195(35);
	sub_wire2(62, 36)    <= sub_wire195(36);
	sub_wire2(62, 37)    <= sub_wire195(37);
	sub_wire2(62, 38)    <= sub_wire195(38);
	sub_wire2(62, 39)    <= sub_wire195(39);
	sub_wire2(61, 0)    <= sub_wire196(0);
	sub_wire2(61, 1)    <= sub_wire196(1);
	sub_wire2(61, 2)    <= sub_wire196(2);
	sub_wire2(61, 3)    <= sub_wire196(3);
	sub_wire2(61, 4)    <= sub_wire196(4);
	sub_wire2(61, 5)    <= sub_wire196(5);
	sub_wire2(61, 6)    <= sub_wire196(6);
	sub_wire2(61, 7)    <= sub_wire196(7);
	sub_wire2(61, 8)    <= sub_wire196(8);
	sub_wire2(61, 9)    <= sub_wire196(9);
	sub_wire2(61, 10)    <= sub_wire196(10);
	sub_wire2(61, 11)    <= sub_wire196(11);
	sub_wire2(61, 12)    <= sub_wire196(12);
	sub_wire2(61, 13)    <= sub_wire196(13);
	sub_wire2(61, 14)    <= sub_wire196(14);
	sub_wire2(61, 15)    <= sub_wire196(15);
	sub_wire2(61, 16)    <= sub_wire196(16);
	sub_wire2(61, 17)    <= sub_wire196(17);
	sub_wire2(61, 18)    <= sub_wire196(18);
	sub_wire2(61, 19)    <= sub_wire196(19);
	sub_wire2(61, 20)    <= sub_wire196(20);
	sub_wire2(61, 21)    <= sub_wire196(21);
	sub_wire2(61, 22)    <= sub_wire196(22);
	sub_wire2(61, 23)    <= sub_wire196(23);
	sub_wire2(61, 24)    <= sub_wire196(24);
	sub_wire2(61, 25)    <= sub_wire196(25);
	sub_wire2(61, 26)    <= sub_wire196(26);
	sub_wire2(61, 27)    <= sub_wire196(27);
	sub_wire2(61, 28)    <= sub_wire196(28);
	sub_wire2(61, 29)    <= sub_wire196(29);
	sub_wire2(61, 30)    <= sub_wire196(30);
	sub_wire2(61, 31)    <= sub_wire196(31);
	sub_wire2(61, 32)    <= sub_wire196(32);
	sub_wire2(61, 33)    <= sub_wire196(33);
	sub_wire2(61, 34)    <= sub_wire196(34);
	sub_wire2(61, 35)    <= sub_wire196(35);
	sub_wire2(61, 36)    <= sub_wire196(36);
	sub_wire2(61, 37)    <= sub_wire196(37);
	sub_wire2(61, 38)    <= sub_wire196(38);
	sub_wire2(61, 39)    <= sub_wire196(39);
	sub_wire2(60, 0)    <= sub_wire197(0);
	sub_wire2(60, 1)    <= sub_wire197(1);
	sub_wire2(60, 2)    <= sub_wire197(2);
	sub_wire2(60, 3)    <= sub_wire197(3);
	sub_wire2(60, 4)    <= sub_wire197(4);
	sub_wire2(60, 5)    <= sub_wire197(5);
	sub_wire2(60, 6)    <= sub_wire197(6);
	sub_wire2(60, 7)    <= sub_wire197(7);
	sub_wire2(60, 8)    <= sub_wire197(8);
	sub_wire2(60, 9)    <= sub_wire197(9);
	sub_wire2(60, 10)    <= sub_wire197(10);
	sub_wire2(60, 11)    <= sub_wire197(11);
	sub_wire2(60, 12)    <= sub_wire197(12);
	sub_wire2(60, 13)    <= sub_wire197(13);
	sub_wire2(60, 14)    <= sub_wire197(14);
	sub_wire2(60, 15)    <= sub_wire197(15);
	sub_wire2(60, 16)    <= sub_wire197(16);
	sub_wire2(60, 17)    <= sub_wire197(17);
	sub_wire2(60, 18)    <= sub_wire197(18);
	sub_wire2(60, 19)    <= sub_wire197(19);
	sub_wire2(60, 20)    <= sub_wire197(20);
	sub_wire2(60, 21)    <= sub_wire197(21);
	sub_wire2(60, 22)    <= sub_wire197(22);
	sub_wire2(60, 23)    <= sub_wire197(23);
	sub_wire2(60, 24)    <= sub_wire197(24);
	sub_wire2(60, 25)    <= sub_wire197(25);
	sub_wire2(60, 26)    <= sub_wire197(26);
	sub_wire2(60, 27)    <= sub_wire197(27);
	sub_wire2(60, 28)    <= sub_wire197(28);
	sub_wire2(60, 29)    <= sub_wire197(29);
	sub_wire2(60, 30)    <= sub_wire197(30);
	sub_wire2(60, 31)    <= sub_wire197(31);
	sub_wire2(60, 32)    <= sub_wire197(32);
	sub_wire2(60, 33)    <= sub_wire197(33);
	sub_wire2(60, 34)    <= sub_wire197(34);
	sub_wire2(60, 35)    <= sub_wire197(35);
	sub_wire2(60, 36)    <= sub_wire197(36);
	sub_wire2(60, 37)    <= sub_wire197(37);
	sub_wire2(60, 38)    <= sub_wire197(38);
	sub_wire2(60, 39)    <= sub_wire197(39);
	sub_wire2(59, 0)    <= sub_wire198(0);
	sub_wire2(59, 1)    <= sub_wire198(1);
	sub_wire2(59, 2)    <= sub_wire198(2);
	sub_wire2(59, 3)    <= sub_wire198(3);
	sub_wire2(59, 4)    <= sub_wire198(4);
	sub_wire2(59, 5)    <= sub_wire198(5);
	sub_wire2(59, 6)    <= sub_wire198(6);
	sub_wire2(59, 7)    <= sub_wire198(7);
	sub_wire2(59, 8)    <= sub_wire198(8);
	sub_wire2(59, 9)    <= sub_wire198(9);
	sub_wire2(59, 10)    <= sub_wire198(10);
	sub_wire2(59, 11)    <= sub_wire198(11);
	sub_wire2(59, 12)    <= sub_wire198(12);
	sub_wire2(59, 13)    <= sub_wire198(13);
	sub_wire2(59, 14)    <= sub_wire198(14);
	sub_wire2(59, 15)    <= sub_wire198(15);
	sub_wire2(59, 16)    <= sub_wire198(16);
	sub_wire2(59, 17)    <= sub_wire198(17);
	sub_wire2(59, 18)    <= sub_wire198(18);
	sub_wire2(59, 19)    <= sub_wire198(19);
	sub_wire2(59, 20)    <= sub_wire198(20);
	sub_wire2(59, 21)    <= sub_wire198(21);
	sub_wire2(59, 22)    <= sub_wire198(22);
	sub_wire2(59, 23)    <= sub_wire198(23);
	sub_wire2(59, 24)    <= sub_wire198(24);
	sub_wire2(59, 25)    <= sub_wire198(25);
	sub_wire2(59, 26)    <= sub_wire198(26);
	sub_wire2(59, 27)    <= sub_wire198(27);
	sub_wire2(59, 28)    <= sub_wire198(28);
	sub_wire2(59, 29)    <= sub_wire198(29);
	sub_wire2(59, 30)    <= sub_wire198(30);
	sub_wire2(59, 31)    <= sub_wire198(31);
	sub_wire2(59, 32)    <= sub_wire198(32);
	sub_wire2(59, 33)    <= sub_wire198(33);
	sub_wire2(59, 34)    <= sub_wire198(34);
	sub_wire2(59, 35)    <= sub_wire198(35);
	sub_wire2(59, 36)    <= sub_wire198(36);
	sub_wire2(59, 37)    <= sub_wire198(37);
	sub_wire2(59, 38)    <= sub_wire198(38);
	sub_wire2(59, 39)    <= sub_wire198(39);
	sub_wire2(58, 0)    <= sub_wire199(0);
	sub_wire2(58, 1)    <= sub_wire199(1);
	sub_wire2(58, 2)    <= sub_wire199(2);
	sub_wire2(58, 3)    <= sub_wire199(3);
	sub_wire2(58, 4)    <= sub_wire199(4);
	sub_wire2(58, 5)    <= sub_wire199(5);
	sub_wire2(58, 6)    <= sub_wire199(6);
	sub_wire2(58, 7)    <= sub_wire199(7);
	sub_wire2(58, 8)    <= sub_wire199(8);
	sub_wire2(58, 9)    <= sub_wire199(9);
	sub_wire2(58, 10)    <= sub_wire199(10);
	sub_wire2(58, 11)    <= sub_wire199(11);
	sub_wire2(58, 12)    <= sub_wire199(12);
	sub_wire2(58, 13)    <= sub_wire199(13);
	sub_wire2(58, 14)    <= sub_wire199(14);
	sub_wire2(58, 15)    <= sub_wire199(15);
	sub_wire2(58, 16)    <= sub_wire199(16);
	sub_wire2(58, 17)    <= sub_wire199(17);
	sub_wire2(58, 18)    <= sub_wire199(18);
	sub_wire2(58, 19)    <= sub_wire199(19);
	sub_wire2(58, 20)    <= sub_wire199(20);
	sub_wire2(58, 21)    <= sub_wire199(21);
	sub_wire2(58, 22)    <= sub_wire199(22);
	sub_wire2(58, 23)    <= sub_wire199(23);
	sub_wire2(58, 24)    <= sub_wire199(24);
	sub_wire2(58, 25)    <= sub_wire199(25);
	sub_wire2(58, 26)    <= sub_wire199(26);
	sub_wire2(58, 27)    <= sub_wire199(27);
	sub_wire2(58, 28)    <= sub_wire199(28);
	sub_wire2(58, 29)    <= sub_wire199(29);
	sub_wire2(58, 30)    <= sub_wire199(30);
	sub_wire2(58, 31)    <= sub_wire199(31);
	sub_wire2(58, 32)    <= sub_wire199(32);
	sub_wire2(58, 33)    <= sub_wire199(33);
	sub_wire2(58, 34)    <= sub_wire199(34);
	sub_wire2(58, 35)    <= sub_wire199(35);
	sub_wire2(58, 36)    <= sub_wire199(36);
	sub_wire2(58, 37)    <= sub_wire199(37);
	sub_wire2(58, 38)    <= sub_wire199(38);
	sub_wire2(58, 39)    <= sub_wire199(39);
	sub_wire2(57, 0)    <= sub_wire200(0);
	sub_wire2(57, 1)    <= sub_wire200(1);
	sub_wire2(57, 2)    <= sub_wire200(2);
	sub_wire2(57, 3)    <= sub_wire200(3);
	sub_wire2(57, 4)    <= sub_wire200(4);
	sub_wire2(57, 5)    <= sub_wire200(5);
	sub_wire2(57, 6)    <= sub_wire200(6);
	sub_wire2(57, 7)    <= sub_wire200(7);
	sub_wire2(57, 8)    <= sub_wire200(8);
	sub_wire2(57, 9)    <= sub_wire200(9);
	sub_wire2(57, 10)    <= sub_wire200(10);
	sub_wire2(57, 11)    <= sub_wire200(11);
	sub_wire2(57, 12)    <= sub_wire200(12);
	sub_wire2(57, 13)    <= sub_wire200(13);
	sub_wire2(57, 14)    <= sub_wire200(14);
	sub_wire2(57, 15)    <= sub_wire200(15);
	sub_wire2(57, 16)    <= sub_wire200(16);
	sub_wire2(57, 17)    <= sub_wire200(17);
	sub_wire2(57, 18)    <= sub_wire200(18);
	sub_wire2(57, 19)    <= sub_wire200(19);
	sub_wire2(57, 20)    <= sub_wire200(20);
	sub_wire2(57, 21)    <= sub_wire200(21);
	sub_wire2(57, 22)    <= sub_wire200(22);
	sub_wire2(57, 23)    <= sub_wire200(23);
	sub_wire2(57, 24)    <= sub_wire200(24);
	sub_wire2(57, 25)    <= sub_wire200(25);
	sub_wire2(57, 26)    <= sub_wire200(26);
	sub_wire2(57, 27)    <= sub_wire200(27);
	sub_wire2(57, 28)    <= sub_wire200(28);
	sub_wire2(57, 29)    <= sub_wire200(29);
	sub_wire2(57, 30)    <= sub_wire200(30);
	sub_wire2(57, 31)    <= sub_wire200(31);
	sub_wire2(57, 32)    <= sub_wire200(32);
	sub_wire2(57, 33)    <= sub_wire200(33);
	sub_wire2(57, 34)    <= sub_wire200(34);
	sub_wire2(57, 35)    <= sub_wire200(35);
	sub_wire2(57, 36)    <= sub_wire200(36);
	sub_wire2(57, 37)    <= sub_wire200(37);
	sub_wire2(57, 38)    <= sub_wire200(38);
	sub_wire2(57, 39)    <= sub_wire200(39);
	sub_wire2(56, 0)    <= sub_wire201(0);
	sub_wire2(56, 1)    <= sub_wire201(1);
	sub_wire2(56, 2)    <= sub_wire201(2);
	sub_wire2(56, 3)    <= sub_wire201(3);
	sub_wire2(56, 4)    <= sub_wire201(4);
	sub_wire2(56, 5)    <= sub_wire201(5);
	sub_wire2(56, 6)    <= sub_wire201(6);
	sub_wire2(56, 7)    <= sub_wire201(7);
	sub_wire2(56, 8)    <= sub_wire201(8);
	sub_wire2(56, 9)    <= sub_wire201(9);
	sub_wire2(56, 10)    <= sub_wire201(10);
	sub_wire2(56, 11)    <= sub_wire201(11);
	sub_wire2(56, 12)    <= sub_wire201(12);
	sub_wire2(56, 13)    <= sub_wire201(13);
	sub_wire2(56, 14)    <= sub_wire201(14);
	sub_wire2(56, 15)    <= sub_wire201(15);
	sub_wire2(56, 16)    <= sub_wire201(16);
	sub_wire2(56, 17)    <= sub_wire201(17);
	sub_wire2(56, 18)    <= sub_wire201(18);
	sub_wire2(56, 19)    <= sub_wire201(19);
	sub_wire2(56, 20)    <= sub_wire201(20);
	sub_wire2(56, 21)    <= sub_wire201(21);
	sub_wire2(56, 22)    <= sub_wire201(22);
	sub_wire2(56, 23)    <= sub_wire201(23);
	sub_wire2(56, 24)    <= sub_wire201(24);
	sub_wire2(56, 25)    <= sub_wire201(25);
	sub_wire2(56, 26)    <= sub_wire201(26);
	sub_wire2(56, 27)    <= sub_wire201(27);
	sub_wire2(56, 28)    <= sub_wire201(28);
	sub_wire2(56, 29)    <= sub_wire201(29);
	sub_wire2(56, 30)    <= sub_wire201(30);
	sub_wire2(56, 31)    <= sub_wire201(31);
	sub_wire2(56, 32)    <= sub_wire201(32);
	sub_wire2(56, 33)    <= sub_wire201(33);
	sub_wire2(56, 34)    <= sub_wire201(34);
	sub_wire2(56, 35)    <= sub_wire201(35);
	sub_wire2(56, 36)    <= sub_wire201(36);
	sub_wire2(56, 37)    <= sub_wire201(37);
	sub_wire2(56, 38)    <= sub_wire201(38);
	sub_wire2(56, 39)    <= sub_wire201(39);
	sub_wire2(55, 0)    <= sub_wire202(0);
	sub_wire2(55, 1)    <= sub_wire202(1);
	sub_wire2(55, 2)    <= sub_wire202(2);
	sub_wire2(55, 3)    <= sub_wire202(3);
	sub_wire2(55, 4)    <= sub_wire202(4);
	sub_wire2(55, 5)    <= sub_wire202(5);
	sub_wire2(55, 6)    <= sub_wire202(6);
	sub_wire2(55, 7)    <= sub_wire202(7);
	sub_wire2(55, 8)    <= sub_wire202(8);
	sub_wire2(55, 9)    <= sub_wire202(9);
	sub_wire2(55, 10)    <= sub_wire202(10);
	sub_wire2(55, 11)    <= sub_wire202(11);
	sub_wire2(55, 12)    <= sub_wire202(12);
	sub_wire2(55, 13)    <= sub_wire202(13);
	sub_wire2(55, 14)    <= sub_wire202(14);
	sub_wire2(55, 15)    <= sub_wire202(15);
	sub_wire2(55, 16)    <= sub_wire202(16);
	sub_wire2(55, 17)    <= sub_wire202(17);
	sub_wire2(55, 18)    <= sub_wire202(18);
	sub_wire2(55, 19)    <= sub_wire202(19);
	sub_wire2(55, 20)    <= sub_wire202(20);
	sub_wire2(55, 21)    <= sub_wire202(21);
	sub_wire2(55, 22)    <= sub_wire202(22);
	sub_wire2(55, 23)    <= sub_wire202(23);
	sub_wire2(55, 24)    <= sub_wire202(24);
	sub_wire2(55, 25)    <= sub_wire202(25);
	sub_wire2(55, 26)    <= sub_wire202(26);
	sub_wire2(55, 27)    <= sub_wire202(27);
	sub_wire2(55, 28)    <= sub_wire202(28);
	sub_wire2(55, 29)    <= sub_wire202(29);
	sub_wire2(55, 30)    <= sub_wire202(30);
	sub_wire2(55, 31)    <= sub_wire202(31);
	sub_wire2(55, 32)    <= sub_wire202(32);
	sub_wire2(55, 33)    <= sub_wire202(33);
	sub_wire2(55, 34)    <= sub_wire202(34);
	sub_wire2(55, 35)    <= sub_wire202(35);
	sub_wire2(55, 36)    <= sub_wire202(36);
	sub_wire2(55, 37)    <= sub_wire202(37);
	sub_wire2(55, 38)    <= sub_wire202(38);
	sub_wire2(55, 39)    <= sub_wire202(39);
	sub_wire2(54, 0)    <= sub_wire203(0);
	sub_wire2(54, 1)    <= sub_wire203(1);
	sub_wire2(54, 2)    <= sub_wire203(2);
	sub_wire2(54, 3)    <= sub_wire203(3);
	sub_wire2(54, 4)    <= sub_wire203(4);
	sub_wire2(54, 5)    <= sub_wire203(5);
	sub_wire2(54, 6)    <= sub_wire203(6);
	sub_wire2(54, 7)    <= sub_wire203(7);
	sub_wire2(54, 8)    <= sub_wire203(8);
	sub_wire2(54, 9)    <= sub_wire203(9);
	sub_wire2(54, 10)    <= sub_wire203(10);
	sub_wire2(54, 11)    <= sub_wire203(11);
	sub_wire2(54, 12)    <= sub_wire203(12);
	sub_wire2(54, 13)    <= sub_wire203(13);
	sub_wire2(54, 14)    <= sub_wire203(14);
	sub_wire2(54, 15)    <= sub_wire203(15);
	sub_wire2(54, 16)    <= sub_wire203(16);
	sub_wire2(54, 17)    <= sub_wire203(17);
	sub_wire2(54, 18)    <= sub_wire203(18);
	sub_wire2(54, 19)    <= sub_wire203(19);
	sub_wire2(54, 20)    <= sub_wire203(20);
	sub_wire2(54, 21)    <= sub_wire203(21);
	sub_wire2(54, 22)    <= sub_wire203(22);
	sub_wire2(54, 23)    <= sub_wire203(23);
	sub_wire2(54, 24)    <= sub_wire203(24);
	sub_wire2(54, 25)    <= sub_wire203(25);
	sub_wire2(54, 26)    <= sub_wire203(26);
	sub_wire2(54, 27)    <= sub_wire203(27);
	sub_wire2(54, 28)    <= sub_wire203(28);
	sub_wire2(54, 29)    <= sub_wire203(29);
	sub_wire2(54, 30)    <= sub_wire203(30);
	sub_wire2(54, 31)    <= sub_wire203(31);
	sub_wire2(54, 32)    <= sub_wire203(32);
	sub_wire2(54, 33)    <= sub_wire203(33);
	sub_wire2(54, 34)    <= sub_wire203(34);
	sub_wire2(54, 35)    <= sub_wire203(35);
	sub_wire2(54, 36)    <= sub_wire203(36);
	sub_wire2(54, 37)    <= sub_wire203(37);
	sub_wire2(54, 38)    <= sub_wire203(38);
	sub_wire2(54, 39)    <= sub_wire203(39);
	sub_wire2(53, 0)    <= sub_wire204(0);
	sub_wire2(53, 1)    <= sub_wire204(1);
	sub_wire2(53, 2)    <= sub_wire204(2);
	sub_wire2(53, 3)    <= sub_wire204(3);
	sub_wire2(53, 4)    <= sub_wire204(4);
	sub_wire2(53, 5)    <= sub_wire204(5);
	sub_wire2(53, 6)    <= sub_wire204(6);
	sub_wire2(53, 7)    <= sub_wire204(7);
	sub_wire2(53, 8)    <= sub_wire204(8);
	sub_wire2(53, 9)    <= sub_wire204(9);
	sub_wire2(53, 10)    <= sub_wire204(10);
	sub_wire2(53, 11)    <= sub_wire204(11);
	sub_wire2(53, 12)    <= sub_wire204(12);
	sub_wire2(53, 13)    <= sub_wire204(13);
	sub_wire2(53, 14)    <= sub_wire204(14);
	sub_wire2(53, 15)    <= sub_wire204(15);
	sub_wire2(53, 16)    <= sub_wire204(16);
	sub_wire2(53, 17)    <= sub_wire204(17);
	sub_wire2(53, 18)    <= sub_wire204(18);
	sub_wire2(53, 19)    <= sub_wire204(19);
	sub_wire2(53, 20)    <= sub_wire204(20);
	sub_wire2(53, 21)    <= sub_wire204(21);
	sub_wire2(53, 22)    <= sub_wire204(22);
	sub_wire2(53, 23)    <= sub_wire204(23);
	sub_wire2(53, 24)    <= sub_wire204(24);
	sub_wire2(53, 25)    <= sub_wire204(25);
	sub_wire2(53, 26)    <= sub_wire204(26);
	sub_wire2(53, 27)    <= sub_wire204(27);
	sub_wire2(53, 28)    <= sub_wire204(28);
	sub_wire2(53, 29)    <= sub_wire204(29);
	sub_wire2(53, 30)    <= sub_wire204(30);
	sub_wire2(53, 31)    <= sub_wire204(31);
	sub_wire2(53, 32)    <= sub_wire204(32);
	sub_wire2(53, 33)    <= sub_wire204(33);
	sub_wire2(53, 34)    <= sub_wire204(34);
	sub_wire2(53, 35)    <= sub_wire204(35);
	sub_wire2(53, 36)    <= sub_wire204(36);
	sub_wire2(53, 37)    <= sub_wire204(37);
	sub_wire2(53, 38)    <= sub_wire204(38);
	sub_wire2(53, 39)    <= sub_wire204(39);
	sub_wire2(52, 0)    <= sub_wire205(0);
	sub_wire2(52, 1)    <= sub_wire205(1);
	sub_wire2(52, 2)    <= sub_wire205(2);
	sub_wire2(52, 3)    <= sub_wire205(3);
	sub_wire2(52, 4)    <= sub_wire205(4);
	sub_wire2(52, 5)    <= sub_wire205(5);
	sub_wire2(52, 6)    <= sub_wire205(6);
	sub_wire2(52, 7)    <= sub_wire205(7);
	sub_wire2(52, 8)    <= sub_wire205(8);
	sub_wire2(52, 9)    <= sub_wire205(9);
	sub_wire2(52, 10)    <= sub_wire205(10);
	sub_wire2(52, 11)    <= sub_wire205(11);
	sub_wire2(52, 12)    <= sub_wire205(12);
	sub_wire2(52, 13)    <= sub_wire205(13);
	sub_wire2(52, 14)    <= sub_wire205(14);
	sub_wire2(52, 15)    <= sub_wire205(15);
	sub_wire2(52, 16)    <= sub_wire205(16);
	sub_wire2(52, 17)    <= sub_wire205(17);
	sub_wire2(52, 18)    <= sub_wire205(18);
	sub_wire2(52, 19)    <= sub_wire205(19);
	sub_wire2(52, 20)    <= sub_wire205(20);
	sub_wire2(52, 21)    <= sub_wire205(21);
	sub_wire2(52, 22)    <= sub_wire205(22);
	sub_wire2(52, 23)    <= sub_wire205(23);
	sub_wire2(52, 24)    <= sub_wire205(24);
	sub_wire2(52, 25)    <= sub_wire205(25);
	sub_wire2(52, 26)    <= sub_wire205(26);
	sub_wire2(52, 27)    <= sub_wire205(27);
	sub_wire2(52, 28)    <= sub_wire205(28);
	sub_wire2(52, 29)    <= sub_wire205(29);
	sub_wire2(52, 30)    <= sub_wire205(30);
	sub_wire2(52, 31)    <= sub_wire205(31);
	sub_wire2(52, 32)    <= sub_wire205(32);
	sub_wire2(52, 33)    <= sub_wire205(33);
	sub_wire2(52, 34)    <= sub_wire205(34);
	sub_wire2(52, 35)    <= sub_wire205(35);
	sub_wire2(52, 36)    <= sub_wire205(36);
	sub_wire2(52, 37)    <= sub_wire205(37);
	sub_wire2(52, 38)    <= sub_wire205(38);
	sub_wire2(52, 39)    <= sub_wire205(39);
	sub_wire2(51, 0)    <= sub_wire206(0);
	sub_wire2(51, 1)    <= sub_wire206(1);
	sub_wire2(51, 2)    <= sub_wire206(2);
	sub_wire2(51, 3)    <= sub_wire206(3);
	sub_wire2(51, 4)    <= sub_wire206(4);
	sub_wire2(51, 5)    <= sub_wire206(5);
	sub_wire2(51, 6)    <= sub_wire206(6);
	sub_wire2(51, 7)    <= sub_wire206(7);
	sub_wire2(51, 8)    <= sub_wire206(8);
	sub_wire2(51, 9)    <= sub_wire206(9);
	sub_wire2(51, 10)    <= sub_wire206(10);
	sub_wire2(51, 11)    <= sub_wire206(11);
	sub_wire2(51, 12)    <= sub_wire206(12);
	sub_wire2(51, 13)    <= sub_wire206(13);
	sub_wire2(51, 14)    <= sub_wire206(14);
	sub_wire2(51, 15)    <= sub_wire206(15);
	sub_wire2(51, 16)    <= sub_wire206(16);
	sub_wire2(51, 17)    <= sub_wire206(17);
	sub_wire2(51, 18)    <= sub_wire206(18);
	sub_wire2(51, 19)    <= sub_wire206(19);
	sub_wire2(51, 20)    <= sub_wire206(20);
	sub_wire2(51, 21)    <= sub_wire206(21);
	sub_wire2(51, 22)    <= sub_wire206(22);
	sub_wire2(51, 23)    <= sub_wire206(23);
	sub_wire2(51, 24)    <= sub_wire206(24);
	sub_wire2(51, 25)    <= sub_wire206(25);
	sub_wire2(51, 26)    <= sub_wire206(26);
	sub_wire2(51, 27)    <= sub_wire206(27);
	sub_wire2(51, 28)    <= sub_wire206(28);
	sub_wire2(51, 29)    <= sub_wire206(29);
	sub_wire2(51, 30)    <= sub_wire206(30);
	sub_wire2(51, 31)    <= sub_wire206(31);
	sub_wire2(51, 32)    <= sub_wire206(32);
	sub_wire2(51, 33)    <= sub_wire206(33);
	sub_wire2(51, 34)    <= sub_wire206(34);
	sub_wire2(51, 35)    <= sub_wire206(35);
	sub_wire2(51, 36)    <= sub_wire206(36);
	sub_wire2(51, 37)    <= sub_wire206(37);
	sub_wire2(51, 38)    <= sub_wire206(38);
	sub_wire2(51, 39)    <= sub_wire206(39);
	sub_wire2(50, 0)    <= sub_wire207(0);
	sub_wire2(50, 1)    <= sub_wire207(1);
	sub_wire2(50, 2)    <= sub_wire207(2);
	sub_wire2(50, 3)    <= sub_wire207(3);
	sub_wire2(50, 4)    <= sub_wire207(4);
	sub_wire2(50, 5)    <= sub_wire207(5);
	sub_wire2(50, 6)    <= sub_wire207(6);
	sub_wire2(50, 7)    <= sub_wire207(7);
	sub_wire2(50, 8)    <= sub_wire207(8);
	sub_wire2(50, 9)    <= sub_wire207(9);
	sub_wire2(50, 10)    <= sub_wire207(10);
	sub_wire2(50, 11)    <= sub_wire207(11);
	sub_wire2(50, 12)    <= sub_wire207(12);
	sub_wire2(50, 13)    <= sub_wire207(13);
	sub_wire2(50, 14)    <= sub_wire207(14);
	sub_wire2(50, 15)    <= sub_wire207(15);
	sub_wire2(50, 16)    <= sub_wire207(16);
	sub_wire2(50, 17)    <= sub_wire207(17);
	sub_wire2(50, 18)    <= sub_wire207(18);
	sub_wire2(50, 19)    <= sub_wire207(19);
	sub_wire2(50, 20)    <= sub_wire207(20);
	sub_wire2(50, 21)    <= sub_wire207(21);
	sub_wire2(50, 22)    <= sub_wire207(22);
	sub_wire2(50, 23)    <= sub_wire207(23);
	sub_wire2(50, 24)    <= sub_wire207(24);
	sub_wire2(50, 25)    <= sub_wire207(25);
	sub_wire2(50, 26)    <= sub_wire207(26);
	sub_wire2(50, 27)    <= sub_wire207(27);
	sub_wire2(50, 28)    <= sub_wire207(28);
	sub_wire2(50, 29)    <= sub_wire207(29);
	sub_wire2(50, 30)    <= sub_wire207(30);
	sub_wire2(50, 31)    <= sub_wire207(31);
	sub_wire2(50, 32)    <= sub_wire207(32);
	sub_wire2(50, 33)    <= sub_wire207(33);
	sub_wire2(50, 34)    <= sub_wire207(34);
	sub_wire2(50, 35)    <= sub_wire207(35);
	sub_wire2(50, 36)    <= sub_wire207(36);
	sub_wire2(50, 37)    <= sub_wire207(37);
	sub_wire2(50, 38)    <= sub_wire207(38);
	sub_wire2(50, 39)    <= sub_wire207(39);
	sub_wire2(49, 0)    <= sub_wire208(0);
	sub_wire2(49, 1)    <= sub_wire208(1);
	sub_wire2(49, 2)    <= sub_wire208(2);
	sub_wire2(49, 3)    <= sub_wire208(3);
	sub_wire2(49, 4)    <= sub_wire208(4);
	sub_wire2(49, 5)    <= sub_wire208(5);
	sub_wire2(49, 6)    <= sub_wire208(6);
	sub_wire2(49, 7)    <= sub_wire208(7);
	sub_wire2(49, 8)    <= sub_wire208(8);
	sub_wire2(49, 9)    <= sub_wire208(9);
	sub_wire2(49, 10)    <= sub_wire208(10);
	sub_wire2(49, 11)    <= sub_wire208(11);
	sub_wire2(49, 12)    <= sub_wire208(12);
	sub_wire2(49, 13)    <= sub_wire208(13);
	sub_wire2(49, 14)    <= sub_wire208(14);
	sub_wire2(49, 15)    <= sub_wire208(15);
	sub_wire2(49, 16)    <= sub_wire208(16);
	sub_wire2(49, 17)    <= sub_wire208(17);
	sub_wire2(49, 18)    <= sub_wire208(18);
	sub_wire2(49, 19)    <= sub_wire208(19);
	sub_wire2(49, 20)    <= sub_wire208(20);
	sub_wire2(49, 21)    <= sub_wire208(21);
	sub_wire2(49, 22)    <= sub_wire208(22);
	sub_wire2(49, 23)    <= sub_wire208(23);
	sub_wire2(49, 24)    <= sub_wire208(24);
	sub_wire2(49, 25)    <= sub_wire208(25);
	sub_wire2(49, 26)    <= sub_wire208(26);
	sub_wire2(49, 27)    <= sub_wire208(27);
	sub_wire2(49, 28)    <= sub_wire208(28);
	sub_wire2(49, 29)    <= sub_wire208(29);
	sub_wire2(49, 30)    <= sub_wire208(30);
	sub_wire2(49, 31)    <= sub_wire208(31);
	sub_wire2(49, 32)    <= sub_wire208(32);
	sub_wire2(49, 33)    <= sub_wire208(33);
	sub_wire2(49, 34)    <= sub_wire208(34);
	sub_wire2(49, 35)    <= sub_wire208(35);
	sub_wire2(49, 36)    <= sub_wire208(36);
	sub_wire2(49, 37)    <= sub_wire208(37);
	sub_wire2(49, 38)    <= sub_wire208(38);
	sub_wire2(49, 39)    <= sub_wire208(39);
	sub_wire2(48, 0)    <= sub_wire209(0);
	sub_wire2(48, 1)    <= sub_wire209(1);
	sub_wire2(48, 2)    <= sub_wire209(2);
	sub_wire2(48, 3)    <= sub_wire209(3);
	sub_wire2(48, 4)    <= sub_wire209(4);
	sub_wire2(48, 5)    <= sub_wire209(5);
	sub_wire2(48, 6)    <= sub_wire209(6);
	sub_wire2(48, 7)    <= sub_wire209(7);
	sub_wire2(48, 8)    <= sub_wire209(8);
	sub_wire2(48, 9)    <= sub_wire209(9);
	sub_wire2(48, 10)    <= sub_wire209(10);
	sub_wire2(48, 11)    <= sub_wire209(11);
	sub_wire2(48, 12)    <= sub_wire209(12);
	sub_wire2(48, 13)    <= sub_wire209(13);
	sub_wire2(48, 14)    <= sub_wire209(14);
	sub_wire2(48, 15)    <= sub_wire209(15);
	sub_wire2(48, 16)    <= sub_wire209(16);
	sub_wire2(48, 17)    <= sub_wire209(17);
	sub_wire2(48, 18)    <= sub_wire209(18);
	sub_wire2(48, 19)    <= sub_wire209(19);
	sub_wire2(48, 20)    <= sub_wire209(20);
	sub_wire2(48, 21)    <= sub_wire209(21);
	sub_wire2(48, 22)    <= sub_wire209(22);
	sub_wire2(48, 23)    <= sub_wire209(23);
	sub_wire2(48, 24)    <= sub_wire209(24);
	sub_wire2(48, 25)    <= sub_wire209(25);
	sub_wire2(48, 26)    <= sub_wire209(26);
	sub_wire2(48, 27)    <= sub_wire209(27);
	sub_wire2(48, 28)    <= sub_wire209(28);
	sub_wire2(48, 29)    <= sub_wire209(29);
	sub_wire2(48, 30)    <= sub_wire209(30);
	sub_wire2(48, 31)    <= sub_wire209(31);
	sub_wire2(48, 32)    <= sub_wire209(32);
	sub_wire2(48, 33)    <= sub_wire209(33);
	sub_wire2(48, 34)    <= sub_wire209(34);
	sub_wire2(48, 35)    <= sub_wire209(35);
	sub_wire2(48, 36)    <= sub_wire209(36);
	sub_wire2(48, 37)    <= sub_wire209(37);
	sub_wire2(48, 38)    <= sub_wire209(38);
	sub_wire2(48, 39)    <= sub_wire209(39);
	sub_wire2(47, 0)    <= sub_wire210(0);
	sub_wire2(47, 1)    <= sub_wire210(1);
	sub_wire2(47, 2)    <= sub_wire210(2);
	sub_wire2(47, 3)    <= sub_wire210(3);
	sub_wire2(47, 4)    <= sub_wire210(4);
	sub_wire2(47, 5)    <= sub_wire210(5);
	sub_wire2(47, 6)    <= sub_wire210(6);
	sub_wire2(47, 7)    <= sub_wire210(7);
	sub_wire2(47, 8)    <= sub_wire210(8);
	sub_wire2(47, 9)    <= sub_wire210(9);
	sub_wire2(47, 10)    <= sub_wire210(10);
	sub_wire2(47, 11)    <= sub_wire210(11);
	sub_wire2(47, 12)    <= sub_wire210(12);
	sub_wire2(47, 13)    <= sub_wire210(13);
	sub_wire2(47, 14)    <= sub_wire210(14);
	sub_wire2(47, 15)    <= sub_wire210(15);
	sub_wire2(47, 16)    <= sub_wire210(16);
	sub_wire2(47, 17)    <= sub_wire210(17);
	sub_wire2(47, 18)    <= sub_wire210(18);
	sub_wire2(47, 19)    <= sub_wire210(19);
	sub_wire2(47, 20)    <= sub_wire210(20);
	sub_wire2(47, 21)    <= sub_wire210(21);
	sub_wire2(47, 22)    <= sub_wire210(22);
	sub_wire2(47, 23)    <= sub_wire210(23);
	sub_wire2(47, 24)    <= sub_wire210(24);
	sub_wire2(47, 25)    <= sub_wire210(25);
	sub_wire2(47, 26)    <= sub_wire210(26);
	sub_wire2(47, 27)    <= sub_wire210(27);
	sub_wire2(47, 28)    <= sub_wire210(28);
	sub_wire2(47, 29)    <= sub_wire210(29);
	sub_wire2(47, 30)    <= sub_wire210(30);
	sub_wire2(47, 31)    <= sub_wire210(31);
	sub_wire2(47, 32)    <= sub_wire210(32);
	sub_wire2(47, 33)    <= sub_wire210(33);
	sub_wire2(47, 34)    <= sub_wire210(34);
	sub_wire2(47, 35)    <= sub_wire210(35);
	sub_wire2(47, 36)    <= sub_wire210(36);
	sub_wire2(47, 37)    <= sub_wire210(37);
	sub_wire2(47, 38)    <= sub_wire210(38);
	sub_wire2(47, 39)    <= sub_wire210(39);
	sub_wire2(46, 0)    <= sub_wire211(0);
	sub_wire2(46, 1)    <= sub_wire211(1);
	sub_wire2(46, 2)    <= sub_wire211(2);
	sub_wire2(46, 3)    <= sub_wire211(3);
	sub_wire2(46, 4)    <= sub_wire211(4);
	sub_wire2(46, 5)    <= sub_wire211(5);
	sub_wire2(46, 6)    <= sub_wire211(6);
	sub_wire2(46, 7)    <= sub_wire211(7);
	sub_wire2(46, 8)    <= sub_wire211(8);
	sub_wire2(46, 9)    <= sub_wire211(9);
	sub_wire2(46, 10)    <= sub_wire211(10);
	sub_wire2(46, 11)    <= sub_wire211(11);
	sub_wire2(46, 12)    <= sub_wire211(12);
	sub_wire2(46, 13)    <= sub_wire211(13);
	sub_wire2(46, 14)    <= sub_wire211(14);
	sub_wire2(46, 15)    <= sub_wire211(15);
	sub_wire2(46, 16)    <= sub_wire211(16);
	sub_wire2(46, 17)    <= sub_wire211(17);
	sub_wire2(46, 18)    <= sub_wire211(18);
	sub_wire2(46, 19)    <= sub_wire211(19);
	sub_wire2(46, 20)    <= sub_wire211(20);
	sub_wire2(46, 21)    <= sub_wire211(21);
	sub_wire2(46, 22)    <= sub_wire211(22);
	sub_wire2(46, 23)    <= sub_wire211(23);
	sub_wire2(46, 24)    <= sub_wire211(24);
	sub_wire2(46, 25)    <= sub_wire211(25);
	sub_wire2(46, 26)    <= sub_wire211(26);
	sub_wire2(46, 27)    <= sub_wire211(27);
	sub_wire2(46, 28)    <= sub_wire211(28);
	sub_wire2(46, 29)    <= sub_wire211(29);
	sub_wire2(46, 30)    <= sub_wire211(30);
	sub_wire2(46, 31)    <= sub_wire211(31);
	sub_wire2(46, 32)    <= sub_wire211(32);
	sub_wire2(46, 33)    <= sub_wire211(33);
	sub_wire2(46, 34)    <= sub_wire211(34);
	sub_wire2(46, 35)    <= sub_wire211(35);
	sub_wire2(46, 36)    <= sub_wire211(36);
	sub_wire2(46, 37)    <= sub_wire211(37);
	sub_wire2(46, 38)    <= sub_wire211(38);
	sub_wire2(46, 39)    <= sub_wire211(39);
	sub_wire2(45, 0)    <= sub_wire212(0);
	sub_wire2(45, 1)    <= sub_wire212(1);
	sub_wire2(45, 2)    <= sub_wire212(2);
	sub_wire2(45, 3)    <= sub_wire212(3);
	sub_wire2(45, 4)    <= sub_wire212(4);
	sub_wire2(45, 5)    <= sub_wire212(5);
	sub_wire2(45, 6)    <= sub_wire212(6);
	sub_wire2(45, 7)    <= sub_wire212(7);
	sub_wire2(45, 8)    <= sub_wire212(8);
	sub_wire2(45, 9)    <= sub_wire212(9);
	sub_wire2(45, 10)    <= sub_wire212(10);
	sub_wire2(45, 11)    <= sub_wire212(11);
	sub_wire2(45, 12)    <= sub_wire212(12);
	sub_wire2(45, 13)    <= sub_wire212(13);
	sub_wire2(45, 14)    <= sub_wire212(14);
	sub_wire2(45, 15)    <= sub_wire212(15);
	sub_wire2(45, 16)    <= sub_wire212(16);
	sub_wire2(45, 17)    <= sub_wire212(17);
	sub_wire2(45, 18)    <= sub_wire212(18);
	sub_wire2(45, 19)    <= sub_wire212(19);
	sub_wire2(45, 20)    <= sub_wire212(20);
	sub_wire2(45, 21)    <= sub_wire212(21);
	sub_wire2(45, 22)    <= sub_wire212(22);
	sub_wire2(45, 23)    <= sub_wire212(23);
	sub_wire2(45, 24)    <= sub_wire212(24);
	sub_wire2(45, 25)    <= sub_wire212(25);
	sub_wire2(45, 26)    <= sub_wire212(26);
	sub_wire2(45, 27)    <= sub_wire212(27);
	sub_wire2(45, 28)    <= sub_wire212(28);
	sub_wire2(45, 29)    <= sub_wire212(29);
	sub_wire2(45, 30)    <= sub_wire212(30);
	sub_wire2(45, 31)    <= sub_wire212(31);
	sub_wire2(45, 32)    <= sub_wire212(32);
	sub_wire2(45, 33)    <= sub_wire212(33);
	sub_wire2(45, 34)    <= sub_wire212(34);
	sub_wire2(45, 35)    <= sub_wire212(35);
	sub_wire2(45, 36)    <= sub_wire212(36);
	sub_wire2(45, 37)    <= sub_wire212(37);
	sub_wire2(45, 38)    <= sub_wire212(38);
	sub_wire2(45, 39)    <= sub_wire212(39);
	sub_wire2(44, 0)    <= sub_wire213(0);
	sub_wire2(44, 1)    <= sub_wire213(1);
	sub_wire2(44, 2)    <= sub_wire213(2);
	sub_wire2(44, 3)    <= sub_wire213(3);
	sub_wire2(44, 4)    <= sub_wire213(4);
	sub_wire2(44, 5)    <= sub_wire213(5);
	sub_wire2(44, 6)    <= sub_wire213(6);
	sub_wire2(44, 7)    <= sub_wire213(7);
	sub_wire2(44, 8)    <= sub_wire213(8);
	sub_wire2(44, 9)    <= sub_wire213(9);
	sub_wire2(44, 10)    <= sub_wire213(10);
	sub_wire2(44, 11)    <= sub_wire213(11);
	sub_wire2(44, 12)    <= sub_wire213(12);
	sub_wire2(44, 13)    <= sub_wire213(13);
	sub_wire2(44, 14)    <= sub_wire213(14);
	sub_wire2(44, 15)    <= sub_wire213(15);
	sub_wire2(44, 16)    <= sub_wire213(16);
	sub_wire2(44, 17)    <= sub_wire213(17);
	sub_wire2(44, 18)    <= sub_wire213(18);
	sub_wire2(44, 19)    <= sub_wire213(19);
	sub_wire2(44, 20)    <= sub_wire213(20);
	sub_wire2(44, 21)    <= sub_wire213(21);
	sub_wire2(44, 22)    <= sub_wire213(22);
	sub_wire2(44, 23)    <= sub_wire213(23);
	sub_wire2(44, 24)    <= sub_wire213(24);
	sub_wire2(44, 25)    <= sub_wire213(25);
	sub_wire2(44, 26)    <= sub_wire213(26);
	sub_wire2(44, 27)    <= sub_wire213(27);
	sub_wire2(44, 28)    <= sub_wire213(28);
	sub_wire2(44, 29)    <= sub_wire213(29);
	sub_wire2(44, 30)    <= sub_wire213(30);
	sub_wire2(44, 31)    <= sub_wire213(31);
	sub_wire2(44, 32)    <= sub_wire213(32);
	sub_wire2(44, 33)    <= sub_wire213(33);
	sub_wire2(44, 34)    <= sub_wire213(34);
	sub_wire2(44, 35)    <= sub_wire213(35);
	sub_wire2(44, 36)    <= sub_wire213(36);
	sub_wire2(44, 37)    <= sub_wire213(37);
	sub_wire2(44, 38)    <= sub_wire213(38);
	sub_wire2(44, 39)    <= sub_wire213(39);
	sub_wire2(43, 0)    <= sub_wire214(0);
	sub_wire2(43, 1)    <= sub_wire214(1);
	sub_wire2(43, 2)    <= sub_wire214(2);
	sub_wire2(43, 3)    <= sub_wire214(3);
	sub_wire2(43, 4)    <= sub_wire214(4);
	sub_wire2(43, 5)    <= sub_wire214(5);
	sub_wire2(43, 6)    <= sub_wire214(6);
	sub_wire2(43, 7)    <= sub_wire214(7);
	sub_wire2(43, 8)    <= sub_wire214(8);
	sub_wire2(43, 9)    <= sub_wire214(9);
	sub_wire2(43, 10)    <= sub_wire214(10);
	sub_wire2(43, 11)    <= sub_wire214(11);
	sub_wire2(43, 12)    <= sub_wire214(12);
	sub_wire2(43, 13)    <= sub_wire214(13);
	sub_wire2(43, 14)    <= sub_wire214(14);
	sub_wire2(43, 15)    <= sub_wire214(15);
	sub_wire2(43, 16)    <= sub_wire214(16);
	sub_wire2(43, 17)    <= sub_wire214(17);
	sub_wire2(43, 18)    <= sub_wire214(18);
	sub_wire2(43, 19)    <= sub_wire214(19);
	sub_wire2(43, 20)    <= sub_wire214(20);
	sub_wire2(43, 21)    <= sub_wire214(21);
	sub_wire2(43, 22)    <= sub_wire214(22);
	sub_wire2(43, 23)    <= sub_wire214(23);
	sub_wire2(43, 24)    <= sub_wire214(24);
	sub_wire2(43, 25)    <= sub_wire214(25);
	sub_wire2(43, 26)    <= sub_wire214(26);
	sub_wire2(43, 27)    <= sub_wire214(27);
	sub_wire2(43, 28)    <= sub_wire214(28);
	sub_wire2(43, 29)    <= sub_wire214(29);
	sub_wire2(43, 30)    <= sub_wire214(30);
	sub_wire2(43, 31)    <= sub_wire214(31);
	sub_wire2(43, 32)    <= sub_wire214(32);
	sub_wire2(43, 33)    <= sub_wire214(33);
	sub_wire2(43, 34)    <= sub_wire214(34);
	sub_wire2(43, 35)    <= sub_wire214(35);
	sub_wire2(43, 36)    <= sub_wire214(36);
	sub_wire2(43, 37)    <= sub_wire214(37);
	sub_wire2(43, 38)    <= sub_wire214(38);
	sub_wire2(43, 39)    <= sub_wire214(39);
	sub_wire2(42, 0)    <= sub_wire215(0);
	sub_wire2(42, 1)    <= sub_wire215(1);
	sub_wire2(42, 2)    <= sub_wire215(2);
	sub_wire2(42, 3)    <= sub_wire215(3);
	sub_wire2(42, 4)    <= sub_wire215(4);
	sub_wire2(42, 5)    <= sub_wire215(5);
	sub_wire2(42, 6)    <= sub_wire215(6);
	sub_wire2(42, 7)    <= sub_wire215(7);
	sub_wire2(42, 8)    <= sub_wire215(8);
	sub_wire2(42, 9)    <= sub_wire215(9);
	sub_wire2(42, 10)    <= sub_wire215(10);
	sub_wire2(42, 11)    <= sub_wire215(11);
	sub_wire2(42, 12)    <= sub_wire215(12);
	sub_wire2(42, 13)    <= sub_wire215(13);
	sub_wire2(42, 14)    <= sub_wire215(14);
	sub_wire2(42, 15)    <= sub_wire215(15);
	sub_wire2(42, 16)    <= sub_wire215(16);
	sub_wire2(42, 17)    <= sub_wire215(17);
	sub_wire2(42, 18)    <= sub_wire215(18);
	sub_wire2(42, 19)    <= sub_wire215(19);
	sub_wire2(42, 20)    <= sub_wire215(20);
	sub_wire2(42, 21)    <= sub_wire215(21);
	sub_wire2(42, 22)    <= sub_wire215(22);
	sub_wire2(42, 23)    <= sub_wire215(23);
	sub_wire2(42, 24)    <= sub_wire215(24);
	sub_wire2(42, 25)    <= sub_wire215(25);
	sub_wire2(42, 26)    <= sub_wire215(26);
	sub_wire2(42, 27)    <= sub_wire215(27);
	sub_wire2(42, 28)    <= sub_wire215(28);
	sub_wire2(42, 29)    <= sub_wire215(29);
	sub_wire2(42, 30)    <= sub_wire215(30);
	sub_wire2(42, 31)    <= sub_wire215(31);
	sub_wire2(42, 32)    <= sub_wire215(32);
	sub_wire2(42, 33)    <= sub_wire215(33);
	sub_wire2(42, 34)    <= sub_wire215(34);
	sub_wire2(42, 35)    <= sub_wire215(35);
	sub_wire2(42, 36)    <= sub_wire215(36);
	sub_wire2(42, 37)    <= sub_wire215(37);
	sub_wire2(42, 38)    <= sub_wire215(38);
	sub_wire2(42, 39)    <= sub_wire215(39);
	sub_wire2(41, 0)    <= sub_wire216(0);
	sub_wire2(41, 1)    <= sub_wire216(1);
	sub_wire2(41, 2)    <= sub_wire216(2);
	sub_wire2(41, 3)    <= sub_wire216(3);
	sub_wire2(41, 4)    <= sub_wire216(4);
	sub_wire2(41, 5)    <= sub_wire216(5);
	sub_wire2(41, 6)    <= sub_wire216(6);
	sub_wire2(41, 7)    <= sub_wire216(7);
	sub_wire2(41, 8)    <= sub_wire216(8);
	sub_wire2(41, 9)    <= sub_wire216(9);
	sub_wire2(41, 10)    <= sub_wire216(10);
	sub_wire2(41, 11)    <= sub_wire216(11);
	sub_wire2(41, 12)    <= sub_wire216(12);
	sub_wire2(41, 13)    <= sub_wire216(13);
	sub_wire2(41, 14)    <= sub_wire216(14);
	sub_wire2(41, 15)    <= sub_wire216(15);
	sub_wire2(41, 16)    <= sub_wire216(16);
	sub_wire2(41, 17)    <= sub_wire216(17);
	sub_wire2(41, 18)    <= sub_wire216(18);
	sub_wire2(41, 19)    <= sub_wire216(19);
	sub_wire2(41, 20)    <= sub_wire216(20);
	sub_wire2(41, 21)    <= sub_wire216(21);
	sub_wire2(41, 22)    <= sub_wire216(22);
	sub_wire2(41, 23)    <= sub_wire216(23);
	sub_wire2(41, 24)    <= sub_wire216(24);
	sub_wire2(41, 25)    <= sub_wire216(25);
	sub_wire2(41, 26)    <= sub_wire216(26);
	sub_wire2(41, 27)    <= sub_wire216(27);
	sub_wire2(41, 28)    <= sub_wire216(28);
	sub_wire2(41, 29)    <= sub_wire216(29);
	sub_wire2(41, 30)    <= sub_wire216(30);
	sub_wire2(41, 31)    <= sub_wire216(31);
	sub_wire2(41, 32)    <= sub_wire216(32);
	sub_wire2(41, 33)    <= sub_wire216(33);
	sub_wire2(41, 34)    <= sub_wire216(34);
	sub_wire2(41, 35)    <= sub_wire216(35);
	sub_wire2(41, 36)    <= sub_wire216(36);
	sub_wire2(41, 37)    <= sub_wire216(37);
	sub_wire2(41, 38)    <= sub_wire216(38);
	sub_wire2(41, 39)    <= sub_wire216(39);
	sub_wire2(40, 0)    <= sub_wire217(0);
	sub_wire2(40, 1)    <= sub_wire217(1);
	sub_wire2(40, 2)    <= sub_wire217(2);
	sub_wire2(40, 3)    <= sub_wire217(3);
	sub_wire2(40, 4)    <= sub_wire217(4);
	sub_wire2(40, 5)    <= sub_wire217(5);
	sub_wire2(40, 6)    <= sub_wire217(6);
	sub_wire2(40, 7)    <= sub_wire217(7);
	sub_wire2(40, 8)    <= sub_wire217(8);
	sub_wire2(40, 9)    <= sub_wire217(9);
	sub_wire2(40, 10)    <= sub_wire217(10);
	sub_wire2(40, 11)    <= sub_wire217(11);
	sub_wire2(40, 12)    <= sub_wire217(12);
	sub_wire2(40, 13)    <= sub_wire217(13);
	sub_wire2(40, 14)    <= sub_wire217(14);
	sub_wire2(40, 15)    <= sub_wire217(15);
	sub_wire2(40, 16)    <= sub_wire217(16);
	sub_wire2(40, 17)    <= sub_wire217(17);
	sub_wire2(40, 18)    <= sub_wire217(18);
	sub_wire2(40, 19)    <= sub_wire217(19);
	sub_wire2(40, 20)    <= sub_wire217(20);
	sub_wire2(40, 21)    <= sub_wire217(21);
	sub_wire2(40, 22)    <= sub_wire217(22);
	sub_wire2(40, 23)    <= sub_wire217(23);
	sub_wire2(40, 24)    <= sub_wire217(24);
	sub_wire2(40, 25)    <= sub_wire217(25);
	sub_wire2(40, 26)    <= sub_wire217(26);
	sub_wire2(40, 27)    <= sub_wire217(27);
	sub_wire2(40, 28)    <= sub_wire217(28);
	sub_wire2(40, 29)    <= sub_wire217(29);
	sub_wire2(40, 30)    <= sub_wire217(30);
	sub_wire2(40, 31)    <= sub_wire217(31);
	sub_wire2(40, 32)    <= sub_wire217(32);
	sub_wire2(40, 33)    <= sub_wire217(33);
	sub_wire2(40, 34)    <= sub_wire217(34);
	sub_wire2(40, 35)    <= sub_wire217(35);
	sub_wire2(40, 36)    <= sub_wire217(36);
	sub_wire2(40, 37)    <= sub_wire217(37);
	sub_wire2(40, 38)    <= sub_wire217(38);
	sub_wire2(40, 39)    <= sub_wire217(39);
	sub_wire2(39, 0)    <= sub_wire218(0);
	sub_wire2(39, 1)    <= sub_wire218(1);
	sub_wire2(39, 2)    <= sub_wire218(2);
	sub_wire2(39, 3)    <= sub_wire218(3);
	sub_wire2(39, 4)    <= sub_wire218(4);
	sub_wire2(39, 5)    <= sub_wire218(5);
	sub_wire2(39, 6)    <= sub_wire218(6);
	sub_wire2(39, 7)    <= sub_wire218(7);
	sub_wire2(39, 8)    <= sub_wire218(8);
	sub_wire2(39, 9)    <= sub_wire218(9);
	sub_wire2(39, 10)    <= sub_wire218(10);
	sub_wire2(39, 11)    <= sub_wire218(11);
	sub_wire2(39, 12)    <= sub_wire218(12);
	sub_wire2(39, 13)    <= sub_wire218(13);
	sub_wire2(39, 14)    <= sub_wire218(14);
	sub_wire2(39, 15)    <= sub_wire218(15);
	sub_wire2(39, 16)    <= sub_wire218(16);
	sub_wire2(39, 17)    <= sub_wire218(17);
	sub_wire2(39, 18)    <= sub_wire218(18);
	sub_wire2(39, 19)    <= sub_wire218(19);
	sub_wire2(39, 20)    <= sub_wire218(20);
	sub_wire2(39, 21)    <= sub_wire218(21);
	sub_wire2(39, 22)    <= sub_wire218(22);
	sub_wire2(39, 23)    <= sub_wire218(23);
	sub_wire2(39, 24)    <= sub_wire218(24);
	sub_wire2(39, 25)    <= sub_wire218(25);
	sub_wire2(39, 26)    <= sub_wire218(26);
	sub_wire2(39, 27)    <= sub_wire218(27);
	sub_wire2(39, 28)    <= sub_wire218(28);
	sub_wire2(39, 29)    <= sub_wire218(29);
	sub_wire2(39, 30)    <= sub_wire218(30);
	sub_wire2(39, 31)    <= sub_wire218(31);
	sub_wire2(39, 32)    <= sub_wire218(32);
	sub_wire2(39, 33)    <= sub_wire218(33);
	sub_wire2(39, 34)    <= sub_wire218(34);
	sub_wire2(39, 35)    <= sub_wire218(35);
	sub_wire2(39, 36)    <= sub_wire218(36);
	sub_wire2(39, 37)    <= sub_wire218(37);
	sub_wire2(39, 38)    <= sub_wire218(38);
	sub_wire2(39, 39)    <= sub_wire218(39);
	sub_wire2(38, 0)    <= sub_wire219(0);
	sub_wire2(38, 1)    <= sub_wire219(1);
	sub_wire2(38, 2)    <= sub_wire219(2);
	sub_wire2(38, 3)    <= sub_wire219(3);
	sub_wire2(38, 4)    <= sub_wire219(4);
	sub_wire2(38, 5)    <= sub_wire219(5);
	sub_wire2(38, 6)    <= sub_wire219(6);
	sub_wire2(38, 7)    <= sub_wire219(7);
	sub_wire2(38, 8)    <= sub_wire219(8);
	sub_wire2(38, 9)    <= sub_wire219(9);
	sub_wire2(38, 10)    <= sub_wire219(10);
	sub_wire2(38, 11)    <= sub_wire219(11);
	sub_wire2(38, 12)    <= sub_wire219(12);
	sub_wire2(38, 13)    <= sub_wire219(13);
	sub_wire2(38, 14)    <= sub_wire219(14);
	sub_wire2(38, 15)    <= sub_wire219(15);
	sub_wire2(38, 16)    <= sub_wire219(16);
	sub_wire2(38, 17)    <= sub_wire219(17);
	sub_wire2(38, 18)    <= sub_wire219(18);
	sub_wire2(38, 19)    <= sub_wire219(19);
	sub_wire2(38, 20)    <= sub_wire219(20);
	sub_wire2(38, 21)    <= sub_wire219(21);
	sub_wire2(38, 22)    <= sub_wire219(22);
	sub_wire2(38, 23)    <= sub_wire219(23);
	sub_wire2(38, 24)    <= sub_wire219(24);
	sub_wire2(38, 25)    <= sub_wire219(25);
	sub_wire2(38, 26)    <= sub_wire219(26);
	sub_wire2(38, 27)    <= sub_wire219(27);
	sub_wire2(38, 28)    <= sub_wire219(28);
	sub_wire2(38, 29)    <= sub_wire219(29);
	sub_wire2(38, 30)    <= sub_wire219(30);
	sub_wire2(38, 31)    <= sub_wire219(31);
	sub_wire2(38, 32)    <= sub_wire219(32);
	sub_wire2(38, 33)    <= sub_wire219(33);
	sub_wire2(38, 34)    <= sub_wire219(34);
	sub_wire2(38, 35)    <= sub_wire219(35);
	sub_wire2(38, 36)    <= sub_wire219(36);
	sub_wire2(38, 37)    <= sub_wire219(37);
	sub_wire2(38, 38)    <= sub_wire219(38);
	sub_wire2(38, 39)    <= sub_wire219(39);
	sub_wire2(37, 0)    <= sub_wire220(0);
	sub_wire2(37, 1)    <= sub_wire220(1);
	sub_wire2(37, 2)    <= sub_wire220(2);
	sub_wire2(37, 3)    <= sub_wire220(3);
	sub_wire2(37, 4)    <= sub_wire220(4);
	sub_wire2(37, 5)    <= sub_wire220(5);
	sub_wire2(37, 6)    <= sub_wire220(6);
	sub_wire2(37, 7)    <= sub_wire220(7);
	sub_wire2(37, 8)    <= sub_wire220(8);
	sub_wire2(37, 9)    <= sub_wire220(9);
	sub_wire2(37, 10)    <= sub_wire220(10);
	sub_wire2(37, 11)    <= sub_wire220(11);
	sub_wire2(37, 12)    <= sub_wire220(12);
	sub_wire2(37, 13)    <= sub_wire220(13);
	sub_wire2(37, 14)    <= sub_wire220(14);
	sub_wire2(37, 15)    <= sub_wire220(15);
	sub_wire2(37, 16)    <= sub_wire220(16);
	sub_wire2(37, 17)    <= sub_wire220(17);
	sub_wire2(37, 18)    <= sub_wire220(18);
	sub_wire2(37, 19)    <= sub_wire220(19);
	sub_wire2(37, 20)    <= sub_wire220(20);
	sub_wire2(37, 21)    <= sub_wire220(21);
	sub_wire2(37, 22)    <= sub_wire220(22);
	sub_wire2(37, 23)    <= sub_wire220(23);
	sub_wire2(37, 24)    <= sub_wire220(24);
	sub_wire2(37, 25)    <= sub_wire220(25);
	sub_wire2(37, 26)    <= sub_wire220(26);
	sub_wire2(37, 27)    <= sub_wire220(27);
	sub_wire2(37, 28)    <= sub_wire220(28);
	sub_wire2(37, 29)    <= sub_wire220(29);
	sub_wire2(37, 30)    <= sub_wire220(30);
	sub_wire2(37, 31)    <= sub_wire220(31);
	sub_wire2(37, 32)    <= sub_wire220(32);
	sub_wire2(37, 33)    <= sub_wire220(33);
	sub_wire2(37, 34)    <= sub_wire220(34);
	sub_wire2(37, 35)    <= sub_wire220(35);
	sub_wire2(37, 36)    <= sub_wire220(36);
	sub_wire2(37, 37)    <= sub_wire220(37);
	sub_wire2(37, 38)    <= sub_wire220(38);
	sub_wire2(37, 39)    <= sub_wire220(39);
	sub_wire2(36, 0)    <= sub_wire221(0);
	sub_wire2(36, 1)    <= sub_wire221(1);
	sub_wire2(36, 2)    <= sub_wire221(2);
	sub_wire2(36, 3)    <= sub_wire221(3);
	sub_wire2(36, 4)    <= sub_wire221(4);
	sub_wire2(36, 5)    <= sub_wire221(5);
	sub_wire2(36, 6)    <= sub_wire221(6);
	sub_wire2(36, 7)    <= sub_wire221(7);
	sub_wire2(36, 8)    <= sub_wire221(8);
	sub_wire2(36, 9)    <= sub_wire221(9);
	sub_wire2(36, 10)    <= sub_wire221(10);
	sub_wire2(36, 11)    <= sub_wire221(11);
	sub_wire2(36, 12)    <= sub_wire221(12);
	sub_wire2(36, 13)    <= sub_wire221(13);
	sub_wire2(36, 14)    <= sub_wire221(14);
	sub_wire2(36, 15)    <= sub_wire221(15);
	sub_wire2(36, 16)    <= sub_wire221(16);
	sub_wire2(36, 17)    <= sub_wire221(17);
	sub_wire2(36, 18)    <= sub_wire221(18);
	sub_wire2(36, 19)    <= sub_wire221(19);
	sub_wire2(36, 20)    <= sub_wire221(20);
	sub_wire2(36, 21)    <= sub_wire221(21);
	sub_wire2(36, 22)    <= sub_wire221(22);
	sub_wire2(36, 23)    <= sub_wire221(23);
	sub_wire2(36, 24)    <= sub_wire221(24);
	sub_wire2(36, 25)    <= sub_wire221(25);
	sub_wire2(36, 26)    <= sub_wire221(26);
	sub_wire2(36, 27)    <= sub_wire221(27);
	sub_wire2(36, 28)    <= sub_wire221(28);
	sub_wire2(36, 29)    <= sub_wire221(29);
	sub_wire2(36, 30)    <= sub_wire221(30);
	sub_wire2(36, 31)    <= sub_wire221(31);
	sub_wire2(36, 32)    <= sub_wire221(32);
	sub_wire2(36, 33)    <= sub_wire221(33);
	sub_wire2(36, 34)    <= sub_wire221(34);
	sub_wire2(36, 35)    <= sub_wire221(35);
	sub_wire2(36, 36)    <= sub_wire221(36);
	sub_wire2(36, 37)    <= sub_wire221(37);
	sub_wire2(36, 38)    <= sub_wire221(38);
	sub_wire2(36, 39)    <= sub_wire221(39);
	sub_wire2(35, 0)    <= sub_wire222(0);
	sub_wire2(35, 1)    <= sub_wire222(1);
	sub_wire2(35, 2)    <= sub_wire222(2);
	sub_wire2(35, 3)    <= sub_wire222(3);
	sub_wire2(35, 4)    <= sub_wire222(4);
	sub_wire2(35, 5)    <= sub_wire222(5);
	sub_wire2(35, 6)    <= sub_wire222(6);
	sub_wire2(35, 7)    <= sub_wire222(7);
	sub_wire2(35, 8)    <= sub_wire222(8);
	sub_wire2(35, 9)    <= sub_wire222(9);
	sub_wire2(35, 10)    <= sub_wire222(10);
	sub_wire2(35, 11)    <= sub_wire222(11);
	sub_wire2(35, 12)    <= sub_wire222(12);
	sub_wire2(35, 13)    <= sub_wire222(13);
	sub_wire2(35, 14)    <= sub_wire222(14);
	sub_wire2(35, 15)    <= sub_wire222(15);
	sub_wire2(35, 16)    <= sub_wire222(16);
	sub_wire2(35, 17)    <= sub_wire222(17);
	sub_wire2(35, 18)    <= sub_wire222(18);
	sub_wire2(35, 19)    <= sub_wire222(19);
	sub_wire2(35, 20)    <= sub_wire222(20);
	sub_wire2(35, 21)    <= sub_wire222(21);
	sub_wire2(35, 22)    <= sub_wire222(22);
	sub_wire2(35, 23)    <= sub_wire222(23);
	sub_wire2(35, 24)    <= sub_wire222(24);
	sub_wire2(35, 25)    <= sub_wire222(25);
	sub_wire2(35, 26)    <= sub_wire222(26);
	sub_wire2(35, 27)    <= sub_wire222(27);
	sub_wire2(35, 28)    <= sub_wire222(28);
	sub_wire2(35, 29)    <= sub_wire222(29);
	sub_wire2(35, 30)    <= sub_wire222(30);
	sub_wire2(35, 31)    <= sub_wire222(31);
	sub_wire2(35, 32)    <= sub_wire222(32);
	sub_wire2(35, 33)    <= sub_wire222(33);
	sub_wire2(35, 34)    <= sub_wire222(34);
	sub_wire2(35, 35)    <= sub_wire222(35);
	sub_wire2(35, 36)    <= sub_wire222(36);
	sub_wire2(35, 37)    <= sub_wire222(37);
	sub_wire2(35, 38)    <= sub_wire222(38);
	sub_wire2(35, 39)    <= sub_wire222(39);
	sub_wire2(34, 0)    <= sub_wire223(0);
	sub_wire2(34, 1)    <= sub_wire223(1);
	sub_wire2(34, 2)    <= sub_wire223(2);
	sub_wire2(34, 3)    <= sub_wire223(3);
	sub_wire2(34, 4)    <= sub_wire223(4);
	sub_wire2(34, 5)    <= sub_wire223(5);
	sub_wire2(34, 6)    <= sub_wire223(6);
	sub_wire2(34, 7)    <= sub_wire223(7);
	sub_wire2(34, 8)    <= sub_wire223(8);
	sub_wire2(34, 9)    <= sub_wire223(9);
	sub_wire2(34, 10)    <= sub_wire223(10);
	sub_wire2(34, 11)    <= sub_wire223(11);
	sub_wire2(34, 12)    <= sub_wire223(12);
	sub_wire2(34, 13)    <= sub_wire223(13);
	sub_wire2(34, 14)    <= sub_wire223(14);
	sub_wire2(34, 15)    <= sub_wire223(15);
	sub_wire2(34, 16)    <= sub_wire223(16);
	sub_wire2(34, 17)    <= sub_wire223(17);
	sub_wire2(34, 18)    <= sub_wire223(18);
	sub_wire2(34, 19)    <= sub_wire223(19);
	sub_wire2(34, 20)    <= sub_wire223(20);
	sub_wire2(34, 21)    <= sub_wire223(21);
	sub_wire2(34, 22)    <= sub_wire223(22);
	sub_wire2(34, 23)    <= sub_wire223(23);
	sub_wire2(34, 24)    <= sub_wire223(24);
	sub_wire2(34, 25)    <= sub_wire223(25);
	sub_wire2(34, 26)    <= sub_wire223(26);
	sub_wire2(34, 27)    <= sub_wire223(27);
	sub_wire2(34, 28)    <= sub_wire223(28);
	sub_wire2(34, 29)    <= sub_wire223(29);
	sub_wire2(34, 30)    <= sub_wire223(30);
	sub_wire2(34, 31)    <= sub_wire223(31);
	sub_wire2(34, 32)    <= sub_wire223(32);
	sub_wire2(34, 33)    <= sub_wire223(33);
	sub_wire2(34, 34)    <= sub_wire223(34);
	sub_wire2(34, 35)    <= sub_wire223(35);
	sub_wire2(34, 36)    <= sub_wire223(36);
	sub_wire2(34, 37)    <= sub_wire223(37);
	sub_wire2(34, 38)    <= sub_wire223(38);
	sub_wire2(34, 39)    <= sub_wire223(39);
	sub_wire2(33, 0)    <= sub_wire224(0);
	sub_wire2(33, 1)    <= sub_wire224(1);
	sub_wire2(33, 2)    <= sub_wire224(2);
	sub_wire2(33, 3)    <= sub_wire224(3);
	sub_wire2(33, 4)    <= sub_wire224(4);
	sub_wire2(33, 5)    <= sub_wire224(5);
	sub_wire2(33, 6)    <= sub_wire224(6);
	sub_wire2(33, 7)    <= sub_wire224(7);
	sub_wire2(33, 8)    <= sub_wire224(8);
	sub_wire2(33, 9)    <= sub_wire224(9);
	sub_wire2(33, 10)    <= sub_wire224(10);
	sub_wire2(33, 11)    <= sub_wire224(11);
	sub_wire2(33, 12)    <= sub_wire224(12);
	sub_wire2(33, 13)    <= sub_wire224(13);
	sub_wire2(33, 14)    <= sub_wire224(14);
	sub_wire2(33, 15)    <= sub_wire224(15);
	sub_wire2(33, 16)    <= sub_wire224(16);
	sub_wire2(33, 17)    <= sub_wire224(17);
	sub_wire2(33, 18)    <= sub_wire224(18);
	sub_wire2(33, 19)    <= sub_wire224(19);
	sub_wire2(33, 20)    <= sub_wire224(20);
	sub_wire2(33, 21)    <= sub_wire224(21);
	sub_wire2(33, 22)    <= sub_wire224(22);
	sub_wire2(33, 23)    <= sub_wire224(23);
	sub_wire2(33, 24)    <= sub_wire224(24);
	sub_wire2(33, 25)    <= sub_wire224(25);
	sub_wire2(33, 26)    <= sub_wire224(26);
	sub_wire2(33, 27)    <= sub_wire224(27);
	sub_wire2(33, 28)    <= sub_wire224(28);
	sub_wire2(33, 29)    <= sub_wire224(29);
	sub_wire2(33, 30)    <= sub_wire224(30);
	sub_wire2(33, 31)    <= sub_wire224(31);
	sub_wire2(33, 32)    <= sub_wire224(32);
	sub_wire2(33, 33)    <= sub_wire224(33);
	sub_wire2(33, 34)    <= sub_wire224(34);
	sub_wire2(33, 35)    <= sub_wire224(35);
	sub_wire2(33, 36)    <= sub_wire224(36);
	sub_wire2(33, 37)    <= sub_wire224(37);
	sub_wire2(33, 38)    <= sub_wire224(38);
	sub_wire2(33, 39)    <= sub_wire224(39);
	sub_wire2(32, 0)    <= sub_wire225(0);
	sub_wire2(32, 1)    <= sub_wire225(1);
	sub_wire2(32, 2)    <= sub_wire225(2);
	sub_wire2(32, 3)    <= sub_wire225(3);
	sub_wire2(32, 4)    <= sub_wire225(4);
	sub_wire2(32, 5)    <= sub_wire225(5);
	sub_wire2(32, 6)    <= sub_wire225(6);
	sub_wire2(32, 7)    <= sub_wire225(7);
	sub_wire2(32, 8)    <= sub_wire225(8);
	sub_wire2(32, 9)    <= sub_wire225(9);
	sub_wire2(32, 10)    <= sub_wire225(10);
	sub_wire2(32, 11)    <= sub_wire225(11);
	sub_wire2(32, 12)    <= sub_wire225(12);
	sub_wire2(32, 13)    <= sub_wire225(13);
	sub_wire2(32, 14)    <= sub_wire225(14);
	sub_wire2(32, 15)    <= sub_wire225(15);
	sub_wire2(32, 16)    <= sub_wire225(16);
	sub_wire2(32, 17)    <= sub_wire225(17);
	sub_wire2(32, 18)    <= sub_wire225(18);
	sub_wire2(32, 19)    <= sub_wire225(19);
	sub_wire2(32, 20)    <= sub_wire225(20);
	sub_wire2(32, 21)    <= sub_wire225(21);
	sub_wire2(32, 22)    <= sub_wire225(22);
	sub_wire2(32, 23)    <= sub_wire225(23);
	sub_wire2(32, 24)    <= sub_wire225(24);
	sub_wire2(32, 25)    <= sub_wire225(25);
	sub_wire2(32, 26)    <= sub_wire225(26);
	sub_wire2(32, 27)    <= sub_wire225(27);
	sub_wire2(32, 28)    <= sub_wire225(28);
	sub_wire2(32, 29)    <= sub_wire225(29);
	sub_wire2(32, 30)    <= sub_wire225(30);
	sub_wire2(32, 31)    <= sub_wire225(31);
	sub_wire2(32, 32)    <= sub_wire225(32);
	sub_wire2(32, 33)    <= sub_wire225(33);
	sub_wire2(32, 34)    <= sub_wire225(34);
	sub_wire2(32, 35)    <= sub_wire225(35);
	sub_wire2(32, 36)    <= sub_wire225(36);
	sub_wire2(32, 37)    <= sub_wire225(37);
	sub_wire2(32, 38)    <= sub_wire225(38);
	sub_wire2(32, 39)    <= sub_wire225(39);
	sub_wire2(31, 0)    <= sub_wire226(0);
	sub_wire2(31, 1)    <= sub_wire226(1);
	sub_wire2(31, 2)    <= sub_wire226(2);
	sub_wire2(31, 3)    <= sub_wire226(3);
	sub_wire2(31, 4)    <= sub_wire226(4);
	sub_wire2(31, 5)    <= sub_wire226(5);
	sub_wire2(31, 6)    <= sub_wire226(6);
	sub_wire2(31, 7)    <= sub_wire226(7);
	sub_wire2(31, 8)    <= sub_wire226(8);
	sub_wire2(31, 9)    <= sub_wire226(9);
	sub_wire2(31, 10)    <= sub_wire226(10);
	sub_wire2(31, 11)    <= sub_wire226(11);
	sub_wire2(31, 12)    <= sub_wire226(12);
	sub_wire2(31, 13)    <= sub_wire226(13);
	sub_wire2(31, 14)    <= sub_wire226(14);
	sub_wire2(31, 15)    <= sub_wire226(15);
	sub_wire2(31, 16)    <= sub_wire226(16);
	sub_wire2(31, 17)    <= sub_wire226(17);
	sub_wire2(31, 18)    <= sub_wire226(18);
	sub_wire2(31, 19)    <= sub_wire226(19);
	sub_wire2(31, 20)    <= sub_wire226(20);
	sub_wire2(31, 21)    <= sub_wire226(21);
	sub_wire2(31, 22)    <= sub_wire226(22);
	sub_wire2(31, 23)    <= sub_wire226(23);
	sub_wire2(31, 24)    <= sub_wire226(24);
	sub_wire2(31, 25)    <= sub_wire226(25);
	sub_wire2(31, 26)    <= sub_wire226(26);
	sub_wire2(31, 27)    <= sub_wire226(27);
	sub_wire2(31, 28)    <= sub_wire226(28);
	sub_wire2(31, 29)    <= sub_wire226(29);
	sub_wire2(31, 30)    <= sub_wire226(30);
	sub_wire2(31, 31)    <= sub_wire226(31);
	sub_wire2(31, 32)    <= sub_wire226(32);
	sub_wire2(31, 33)    <= sub_wire226(33);
	sub_wire2(31, 34)    <= sub_wire226(34);
	sub_wire2(31, 35)    <= sub_wire226(35);
	sub_wire2(31, 36)    <= sub_wire226(36);
	sub_wire2(31, 37)    <= sub_wire226(37);
	sub_wire2(31, 38)    <= sub_wire226(38);
	sub_wire2(31, 39)    <= sub_wire226(39);
	sub_wire2(30, 0)    <= sub_wire227(0);
	sub_wire2(30, 1)    <= sub_wire227(1);
	sub_wire2(30, 2)    <= sub_wire227(2);
	sub_wire2(30, 3)    <= sub_wire227(3);
	sub_wire2(30, 4)    <= sub_wire227(4);
	sub_wire2(30, 5)    <= sub_wire227(5);
	sub_wire2(30, 6)    <= sub_wire227(6);
	sub_wire2(30, 7)    <= sub_wire227(7);
	sub_wire2(30, 8)    <= sub_wire227(8);
	sub_wire2(30, 9)    <= sub_wire227(9);
	sub_wire2(30, 10)    <= sub_wire227(10);
	sub_wire2(30, 11)    <= sub_wire227(11);
	sub_wire2(30, 12)    <= sub_wire227(12);
	sub_wire2(30, 13)    <= sub_wire227(13);
	sub_wire2(30, 14)    <= sub_wire227(14);
	sub_wire2(30, 15)    <= sub_wire227(15);
	sub_wire2(30, 16)    <= sub_wire227(16);
	sub_wire2(30, 17)    <= sub_wire227(17);
	sub_wire2(30, 18)    <= sub_wire227(18);
	sub_wire2(30, 19)    <= sub_wire227(19);
	sub_wire2(30, 20)    <= sub_wire227(20);
	sub_wire2(30, 21)    <= sub_wire227(21);
	sub_wire2(30, 22)    <= sub_wire227(22);
	sub_wire2(30, 23)    <= sub_wire227(23);
	sub_wire2(30, 24)    <= sub_wire227(24);
	sub_wire2(30, 25)    <= sub_wire227(25);
	sub_wire2(30, 26)    <= sub_wire227(26);
	sub_wire2(30, 27)    <= sub_wire227(27);
	sub_wire2(30, 28)    <= sub_wire227(28);
	sub_wire2(30, 29)    <= sub_wire227(29);
	sub_wire2(30, 30)    <= sub_wire227(30);
	sub_wire2(30, 31)    <= sub_wire227(31);
	sub_wire2(30, 32)    <= sub_wire227(32);
	sub_wire2(30, 33)    <= sub_wire227(33);
	sub_wire2(30, 34)    <= sub_wire227(34);
	sub_wire2(30, 35)    <= sub_wire227(35);
	sub_wire2(30, 36)    <= sub_wire227(36);
	sub_wire2(30, 37)    <= sub_wire227(37);
	sub_wire2(30, 38)    <= sub_wire227(38);
	sub_wire2(30, 39)    <= sub_wire227(39);
	sub_wire2(29, 0)    <= sub_wire228(0);
	sub_wire2(29, 1)    <= sub_wire228(1);
	sub_wire2(29, 2)    <= sub_wire228(2);
	sub_wire2(29, 3)    <= sub_wire228(3);
	sub_wire2(29, 4)    <= sub_wire228(4);
	sub_wire2(29, 5)    <= sub_wire228(5);
	sub_wire2(29, 6)    <= sub_wire228(6);
	sub_wire2(29, 7)    <= sub_wire228(7);
	sub_wire2(29, 8)    <= sub_wire228(8);
	sub_wire2(29, 9)    <= sub_wire228(9);
	sub_wire2(29, 10)    <= sub_wire228(10);
	sub_wire2(29, 11)    <= sub_wire228(11);
	sub_wire2(29, 12)    <= sub_wire228(12);
	sub_wire2(29, 13)    <= sub_wire228(13);
	sub_wire2(29, 14)    <= sub_wire228(14);
	sub_wire2(29, 15)    <= sub_wire228(15);
	sub_wire2(29, 16)    <= sub_wire228(16);
	sub_wire2(29, 17)    <= sub_wire228(17);
	sub_wire2(29, 18)    <= sub_wire228(18);
	sub_wire2(29, 19)    <= sub_wire228(19);
	sub_wire2(29, 20)    <= sub_wire228(20);
	sub_wire2(29, 21)    <= sub_wire228(21);
	sub_wire2(29, 22)    <= sub_wire228(22);
	sub_wire2(29, 23)    <= sub_wire228(23);
	sub_wire2(29, 24)    <= sub_wire228(24);
	sub_wire2(29, 25)    <= sub_wire228(25);
	sub_wire2(29, 26)    <= sub_wire228(26);
	sub_wire2(29, 27)    <= sub_wire228(27);
	sub_wire2(29, 28)    <= sub_wire228(28);
	sub_wire2(29, 29)    <= sub_wire228(29);
	sub_wire2(29, 30)    <= sub_wire228(30);
	sub_wire2(29, 31)    <= sub_wire228(31);
	sub_wire2(29, 32)    <= sub_wire228(32);
	sub_wire2(29, 33)    <= sub_wire228(33);
	sub_wire2(29, 34)    <= sub_wire228(34);
	sub_wire2(29, 35)    <= sub_wire228(35);
	sub_wire2(29, 36)    <= sub_wire228(36);
	sub_wire2(29, 37)    <= sub_wire228(37);
	sub_wire2(29, 38)    <= sub_wire228(38);
	sub_wire2(29, 39)    <= sub_wire228(39);
	sub_wire2(28, 0)    <= sub_wire229(0);
	sub_wire2(28, 1)    <= sub_wire229(1);
	sub_wire2(28, 2)    <= sub_wire229(2);
	sub_wire2(28, 3)    <= sub_wire229(3);
	sub_wire2(28, 4)    <= sub_wire229(4);
	sub_wire2(28, 5)    <= sub_wire229(5);
	sub_wire2(28, 6)    <= sub_wire229(6);
	sub_wire2(28, 7)    <= sub_wire229(7);
	sub_wire2(28, 8)    <= sub_wire229(8);
	sub_wire2(28, 9)    <= sub_wire229(9);
	sub_wire2(28, 10)    <= sub_wire229(10);
	sub_wire2(28, 11)    <= sub_wire229(11);
	sub_wire2(28, 12)    <= sub_wire229(12);
	sub_wire2(28, 13)    <= sub_wire229(13);
	sub_wire2(28, 14)    <= sub_wire229(14);
	sub_wire2(28, 15)    <= sub_wire229(15);
	sub_wire2(28, 16)    <= sub_wire229(16);
	sub_wire2(28, 17)    <= sub_wire229(17);
	sub_wire2(28, 18)    <= sub_wire229(18);
	sub_wire2(28, 19)    <= sub_wire229(19);
	sub_wire2(28, 20)    <= sub_wire229(20);
	sub_wire2(28, 21)    <= sub_wire229(21);
	sub_wire2(28, 22)    <= sub_wire229(22);
	sub_wire2(28, 23)    <= sub_wire229(23);
	sub_wire2(28, 24)    <= sub_wire229(24);
	sub_wire2(28, 25)    <= sub_wire229(25);
	sub_wire2(28, 26)    <= sub_wire229(26);
	sub_wire2(28, 27)    <= sub_wire229(27);
	sub_wire2(28, 28)    <= sub_wire229(28);
	sub_wire2(28, 29)    <= sub_wire229(29);
	sub_wire2(28, 30)    <= sub_wire229(30);
	sub_wire2(28, 31)    <= sub_wire229(31);
	sub_wire2(28, 32)    <= sub_wire229(32);
	sub_wire2(28, 33)    <= sub_wire229(33);
	sub_wire2(28, 34)    <= sub_wire229(34);
	sub_wire2(28, 35)    <= sub_wire229(35);
	sub_wire2(28, 36)    <= sub_wire229(36);
	sub_wire2(28, 37)    <= sub_wire229(37);
	sub_wire2(28, 38)    <= sub_wire229(38);
	sub_wire2(28, 39)    <= sub_wire229(39);
	sub_wire2(27, 0)    <= sub_wire230(0);
	sub_wire2(27, 1)    <= sub_wire230(1);
	sub_wire2(27, 2)    <= sub_wire230(2);
	sub_wire2(27, 3)    <= sub_wire230(3);
	sub_wire2(27, 4)    <= sub_wire230(4);
	sub_wire2(27, 5)    <= sub_wire230(5);
	sub_wire2(27, 6)    <= sub_wire230(6);
	sub_wire2(27, 7)    <= sub_wire230(7);
	sub_wire2(27, 8)    <= sub_wire230(8);
	sub_wire2(27, 9)    <= sub_wire230(9);
	sub_wire2(27, 10)    <= sub_wire230(10);
	sub_wire2(27, 11)    <= sub_wire230(11);
	sub_wire2(27, 12)    <= sub_wire230(12);
	sub_wire2(27, 13)    <= sub_wire230(13);
	sub_wire2(27, 14)    <= sub_wire230(14);
	sub_wire2(27, 15)    <= sub_wire230(15);
	sub_wire2(27, 16)    <= sub_wire230(16);
	sub_wire2(27, 17)    <= sub_wire230(17);
	sub_wire2(27, 18)    <= sub_wire230(18);
	sub_wire2(27, 19)    <= sub_wire230(19);
	sub_wire2(27, 20)    <= sub_wire230(20);
	sub_wire2(27, 21)    <= sub_wire230(21);
	sub_wire2(27, 22)    <= sub_wire230(22);
	sub_wire2(27, 23)    <= sub_wire230(23);
	sub_wire2(27, 24)    <= sub_wire230(24);
	sub_wire2(27, 25)    <= sub_wire230(25);
	sub_wire2(27, 26)    <= sub_wire230(26);
	sub_wire2(27, 27)    <= sub_wire230(27);
	sub_wire2(27, 28)    <= sub_wire230(28);
	sub_wire2(27, 29)    <= sub_wire230(29);
	sub_wire2(27, 30)    <= sub_wire230(30);
	sub_wire2(27, 31)    <= sub_wire230(31);
	sub_wire2(27, 32)    <= sub_wire230(32);
	sub_wire2(27, 33)    <= sub_wire230(33);
	sub_wire2(27, 34)    <= sub_wire230(34);
	sub_wire2(27, 35)    <= sub_wire230(35);
	sub_wire2(27, 36)    <= sub_wire230(36);
	sub_wire2(27, 37)    <= sub_wire230(37);
	sub_wire2(27, 38)    <= sub_wire230(38);
	sub_wire2(27, 39)    <= sub_wire230(39);
	sub_wire2(26, 0)    <= sub_wire231(0);
	sub_wire2(26, 1)    <= sub_wire231(1);
	sub_wire2(26, 2)    <= sub_wire231(2);
	sub_wire2(26, 3)    <= sub_wire231(3);
	sub_wire2(26, 4)    <= sub_wire231(4);
	sub_wire2(26, 5)    <= sub_wire231(5);
	sub_wire2(26, 6)    <= sub_wire231(6);
	sub_wire2(26, 7)    <= sub_wire231(7);
	sub_wire2(26, 8)    <= sub_wire231(8);
	sub_wire2(26, 9)    <= sub_wire231(9);
	sub_wire2(26, 10)    <= sub_wire231(10);
	sub_wire2(26, 11)    <= sub_wire231(11);
	sub_wire2(26, 12)    <= sub_wire231(12);
	sub_wire2(26, 13)    <= sub_wire231(13);
	sub_wire2(26, 14)    <= sub_wire231(14);
	sub_wire2(26, 15)    <= sub_wire231(15);
	sub_wire2(26, 16)    <= sub_wire231(16);
	sub_wire2(26, 17)    <= sub_wire231(17);
	sub_wire2(26, 18)    <= sub_wire231(18);
	sub_wire2(26, 19)    <= sub_wire231(19);
	sub_wire2(26, 20)    <= sub_wire231(20);
	sub_wire2(26, 21)    <= sub_wire231(21);
	sub_wire2(26, 22)    <= sub_wire231(22);
	sub_wire2(26, 23)    <= sub_wire231(23);
	sub_wire2(26, 24)    <= sub_wire231(24);
	sub_wire2(26, 25)    <= sub_wire231(25);
	sub_wire2(26, 26)    <= sub_wire231(26);
	sub_wire2(26, 27)    <= sub_wire231(27);
	sub_wire2(26, 28)    <= sub_wire231(28);
	sub_wire2(26, 29)    <= sub_wire231(29);
	sub_wire2(26, 30)    <= sub_wire231(30);
	sub_wire2(26, 31)    <= sub_wire231(31);
	sub_wire2(26, 32)    <= sub_wire231(32);
	sub_wire2(26, 33)    <= sub_wire231(33);
	sub_wire2(26, 34)    <= sub_wire231(34);
	sub_wire2(26, 35)    <= sub_wire231(35);
	sub_wire2(26, 36)    <= sub_wire231(36);
	sub_wire2(26, 37)    <= sub_wire231(37);
	sub_wire2(26, 38)    <= sub_wire231(38);
	sub_wire2(26, 39)    <= sub_wire231(39);
	sub_wire2(25, 0)    <= sub_wire232(0);
	sub_wire2(25, 1)    <= sub_wire232(1);
	sub_wire2(25, 2)    <= sub_wire232(2);
	sub_wire2(25, 3)    <= sub_wire232(3);
	sub_wire2(25, 4)    <= sub_wire232(4);
	sub_wire2(25, 5)    <= sub_wire232(5);
	sub_wire2(25, 6)    <= sub_wire232(6);
	sub_wire2(25, 7)    <= sub_wire232(7);
	sub_wire2(25, 8)    <= sub_wire232(8);
	sub_wire2(25, 9)    <= sub_wire232(9);
	sub_wire2(25, 10)    <= sub_wire232(10);
	sub_wire2(25, 11)    <= sub_wire232(11);
	sub_wire2(25, 12)    <= sub_wire232(12);
	sub_wire2(25, 13)    <= sub_wire232(13);
	sub_wire2(25, 14)    <= sub_wire232(14);
	sub_wire2(25, 15)    <= sub_wire232(15);
	sub_wire2(25, 16)    <= sub_wire232(16);
	sub_wire2(25, 17)    <= sub_wire232(17);
	sub_wire2(25, 18)    <= sub_wire232(18);
	sub_wire2(25, 19)    <= sub_wire232(19);
	sub_wire2(25, 20)    <= sub_wire232(20);
	sub_wire2(25, 21)    <= sub_wire232(21);
	sub_wire2(25, 22)    <= sub_wire232(22);
	sub_wire2(25, 23)    <= sub_wire232(23);
	sub_wire2(25, 24)    <= sub_wire232(24);
	sub_wire2(25, 25)    <= sub_wire232(25);
	sub_wire2(25, 26)    <= sub_wire232(26);
	sub_wire2(25, 27)    <= sub_wire232(27);
	sub_wire2(25, 28)    <= sub_wire232(28);
	sub_wire2(25, 29)    <= sub_wire232(29);
	sub_wire2(25, 30)    <= sub_wire232(30);
	sub_wire2(25, 31)    <= sub_wire232(31);
	sub_wire2(25, 32)    <= sub_wire232(32);
	sub_wire2(25, 33)    <= sub_wire232(33);
	sub_wire2(25, 34)    <= sub_wire232(34);
	sub_wire2(25, 35)    <= sub_wire232(35);
	sub_wire2(25, 36)    <= sub_wire232(36);
	sub_wire2(25, 37)    <= sub_wire232(37);
	sub_wire2(25, 38)    <= sub_wire232(38);
	sub_wire2(25, 39)    <= sub_wire232(39);
	sub_wire2(24, 0)    <= sub_wire233(0);
	sub_wire2(24, 1)    <= sub_wire233(1);
	sub_wire2(24, 2)    <= sub_wire233(2);
	sub_wire2(24, 3)    <= sub_wire233(3);
	sub_wire2(24, 4)    <= sub_wire233(4);
	sub_wire2(24, 5)    <= sub_wire233(5);
	sub_wire2(24, 6)    <= sub_wire233(6);
	sub_wire2(24, 7)    <= sub_wire233(7);
	sub_wire2(24, 8)    <= sub_wire233(8);
	sub_wire2(24, 9)    <= sub_wire233(9);
	sub_wire2(24, 10)    <= sub_wire233(10);
	sub_wire2(24, 11)    <= sub_wire233(11);
	sub_wire2(24, 12)    <= sub_wire233(12);
	sub_wire2(24, 13)    <= sub_wire233(13);
	sub_wire2(24, 14)    <= sub_wire233(14);
	sub_wire2(24, 15)    <= sub_wire233(15);
	sub_wire2(24, 16)    <= sub_wire233(16);
	sub_wire2(24, 17)    <= sub_wire233(17);
	sub_wire2(24, 18)    <= sub_wire233(18);
	sub_wire2(24, 19)    <= sub_wire233(19);
	sub_wire2(24, 20)    <= sub_wire233(20);
	sub_wire2(24, 21)    <= sub_wire233(21);
	sub_wire2(24, 22)    <= sub_wire233(22);
	sub_wire2(24, 23)    <= sub_wire233(23);
	sub_wire2(24, 24)    <= sub_wire233(24);
	sub_wire2(24, 25)    <= sub_wire233(25);
	sub_wire2(24, 26)    <= sub_wire233(26);
	sub_wire2(24, 27)    <= sub_wire233(27);
	sub_wire2(24, 28)    <= sub_wire233(28);
	sub_wire2(24, 29)    <= sub_wire233(29);
	sub_wire2(24, 30)    <= sub_wire233(30);
	sub_wire2(24, 31)    <= sub_wire233(31);
	sub_wire2(24, 32)    <= sub_wire233(32);
	sub_wire2(24, 33)    <= sub_wire233(33);
	sub_wire2(24, 34)    <= sub_wire233(34);
	sub_wire2(24, 35)    <= sub_wire233(35);
	sub_wire2(24, 36)    <= sub_wire233(36);
	sub_wire2(24, 37)    <= sub_wire233(37);
	sub_wire2(24, 38)    <= sub_wire233(38);
	sub_wire2(24, 39)    <= sub_wire233(39);
	sub_wire2(23, 0)    <= sub_wire234(0);
	sub_wire2(23, 1)    <= sub_wire234(1);
	sub_wire2(23, 2)    <= sub_wire234(2);
	sub_wire2(23, 3)    <= sub_wire234(3);
	sub_wire2(23, 4)    <= sub_wire234(4);
	sub_wire2(23, 5)    <= sub_wire234(5);
	sub_wire2(23, 6)    <= sub_wire234(6);
	sub_wire2(23, 7)    <= sub_wire234(7);
	sub_wire2(23, 8)    <= sub_wire234(8);
	sub_wire2(23, 9)    <= sub_wire234(9);
	sub_wire2(23, 10)    <= sub_wire234(10);
	sub_wire2(23, 11)    <= sub_wire234(11);
	sub_wire2(23, 12)    <= sub_wire234(12);
	sub_wire2(23, 13)    <= sub_wire234(13);
	sub_wire2(23, 14)    <= sub_wire234(14);
	sub_wire2(23, 15)    <= sub_wire234(15);
	sub_wire2(23, 16)    <= sub_wire234(16);
	sub_wire2(23, 17)    <= sub_wire234(17);
	sub_wire2(23, 18)    <= sub_wire234(18);
	sub_wire2(23, 19)    <= sub_wire234(19);
	sub_wire2(23, 20)    <= sub_wire234(20);
	sub_wire2(23, 21)    <= sub_wire234(21);
	sub_wire2(23, 22)    <= sub_wire234(22);
	sub_wire2(23, 23)    <= sub_wire234(23);
	sub_wire2(23, 24)    <= sub_wire234(24);
	sub_wire2(23, 25)    <= sub_wire234(25);
	sub_wire2(23, 26)    <= sub_wire234(26);
	sub_wire2(23, 27)    <= sub_wire234(27);
	sub_wire2(23, 28)    <= sub_wire234(28);
	sub_wire2(23, 29)    <= sub_wire234(29);
	sub_wire2(23, 30)    <= sub_wire234(30);
	sub_wire2(23, 31)    <= sub_wire234(31);
	sub_wire2(23, 32)    <= sub_wire234(32);
	sub_wire2(23, 33)    <= sub_wire234(33);
	sub_wire2(23, 34)    <= sub_wire234(34);
	sub_wire2(23, 35)    <= sub_wire234(35);
	sub_wire2(23, 36)    <= sub_wire234(36);
	sub_wire2(23, 37)    <= sub_wire234(37);
	sub_wire2(23, 38)    <= sub_wire234(38);
	sub_wire2(23, 39)    <= sub_wire234(39);
	sub_wire2(22, 0)    <= sub_wire235(0);
	sub_wire2(22, 1)    <= sub_wire235(1);
	sub_wire2(22, 2)    <= sub_wire235(2);
	sub_wire2(22, 3)    <= sub_wire235(3);
	sub_wire2(22, 4)    <= sub_wire235(4);
	sub_wire2(22, 5)    <= sub_wire235(5);
	sub_wire2(22, 6)    <= sub_wire235(6);
	sub_wire2(22, 7)    <= sub_wire235(7);
	sub_wire2(22, 8)    <= sub_wire235(8);
	sub_wire2(22, 9)    <= sub_wire235(9);
	sub_wire2(22, 10)    <= sub_wire235(10);
	sub_wire2(22, 11)    <= sub_wire235(11);
	sub_wire2(22, 12)    <= sub_wire235(12);
	sub_wire2(22, 13)    <= sub_wire235(13);
	sub_wire2(22, 14)    <= sub_wire235(14);
	sub_wire2(22, 15)    <= sub_wire235(15);
	sub_wire2(22, 16)    <= sub_wire235(16);
	sub_wire2(22, 17)    <= sub_wire235(17);
	sub_wire2(22, 18)    <= sub_wire235(18);
	sub_wire2(22, 19)    <= sub_wire235(19);
	sub_wire2(22, 20)    <= sub_wire235(20);
	sub_wire2(22, 21)    <= sub_wire235(21);
	sub_wire2(22, 22)    <= sub_wire235(22);
	sub_wire2(22, 23)    <= sub_wire235(23);
	sub_wire2(22, 24)    <= sub_wire235(24);
	sub_wire2(22, 25)    <= sub_wire235(25);
	sub_wire2(22, 26)    <= sub_wire235(26);
	sub_wire2(22, 27)    <= sub_wire235(27);
	sub_wire2(22, 28)    <= sub_wire235(28);
	sub_wire2(22, 29)    <= sub_wire235(29);
	sub_wire2(22, 30)    <= sub_wire235(30);
	sub_wire2(22, 31)    <= sub_wire235(31);
	sub_wire2(22, 32)    <= sub_wire235(32);
	sub_wire2(22, 33)    <= sub_wire235(33);
	sub_wire2(22, 34)    <= sub_wire235(34);
	sub_wire2(22, 35)    <= sub_wire235(35);
	sub_wire2(22, 36)    <= sub_wire235(36);
	sub_wire2(22, 37)    <= sub_wire235(37);
	sub_wire2(22, 38)    <= sub_wire235(38);
	sub_wire2(22, 39)    <= sub_wire235(39);
	sub_wire2(21, 0)    <= sub_wire236(0);
	sub_wire2(21, 1)    <= sub_wire236(1);
	sub_wire2(21, 2)    <= sub_wire236(2);
	sub_wire2(21, 3)    <= sub_wire236(3);
	sub_wire2(21, 4)    <= sub_wire236(4);
	sub_wire2(21, 5)    <= sub_wire236(5);
	sub_wire2(21, 6)    <= sub_wire236(6);
	sub_wire2(21, 7)    <= sub_wire236(7);
	sub_wire2(21, 8)    <= sub_wire236(8);
	sub_wire2(21, 9)    <= sub_wire236(9);
	sub_wire2(21, 10)    <= sub_wire236(10);
	sub_wire2(21, 11)    <= sub_wire236(11);
	sub_wire2(21, 12)    <= sub_wire236(12);
	sub_wire2(21, 13)    <= sub_wire236(13);
	sub_wire2(21, 14)    <= sub_wire236(14);
	sub_wire2(21, 15)    <= sub_wire236(15);
	sub_wire2(21, 16)    <= sub_wire236(16);
	sub_wire2(21, 17)    <= sub_wire236(17);
	sub_wire2(21, 18)    <= sub_wire236(18);
	sub_wire2(21, 19)    <= sub_wire236(19);
	sub_wire2(21, 20)    <= sub_wire236(20);
	sub_wire2(21, 21)    <= sub_wire236(21);
	sub_wire2(21, 22)    <= sub_wire236(22);
	sub_wire2(21, 23)    <= sub_wire236(23);
	sub_wire2(21, 24)    <= sub_wire236(24);
	sub_wire2(21, 25)    <= sub_wire236(25);
	sub_wire2(21, 26)    <= sub_wire236(26);
	sub_wire2(21, 27)    <= sub_wire236(27);
	sub_wire2(21, 28)    <= sub_wire236(28);
	sub_wire2(21, 29)    <= sub_wire236(29);
	sub_wire2(21, 30)    <= sub_wire236(30);
	sub_wire2(21, 31)    <= sub_wire236(31);
	sub_wire2(21, 32)    <= sub_wire236(32);
	sub_wire2(21, 33)    <= sub_wire236(33);
	sub_wire2(21, 34)    <= sub_wire236(34);
	sub_wire2(21, 35)    <= sub_wire236(35);
	sub_wire2(21, 36)    <= sub_wire236(36);
	sub_wire2(21, 37)    <= sub_wire236(37);
	sub_wire2(21, 38)    <= sub_wire236(38);
	sub_wire2(21, 39)    <= sub_wire236(39);
	sub_wire2(20, 0)    <= sub_wire237(0);
	sub_wire2(20, 1)    <= sub_wire237(1);
	sub_wire2(20, 2)    <= sub_wire237(2);
	sub_wire2(20, 3)    <= sub_wire237(3);
	sub_wire2(20, 4)    <= sub_wire237(4);
	sub_wire2(20, 5)    <= sub_wire237(5);
	sub_wire2(20, 6)    <= sub_wire237(6);
	sub_wire2(20, 7)    <= sub_wire237(7);
	sub_wire2(20, 8)    <= sub_wire237(8);
	sub_wire2(20, 9)    <= sub_wire237(9);
	sub_wire2(20, 10)    <= sub_wire237(10);
	sub_wire2(20, 11)    <= sub_wire237(11);
	sub_wire2(20, 12)    <= sub_wire237(12);
	sub_wire2(20, 13)    <= sub_wire237(13);
	sub_wire2(20, 14)    <= sub_wire237(14);
	sub_wire2(20, 15)    <= sub_wire237(15);
	sub_wire2(20, 16)    <= sub_wire237(16);
	sub_wire2(20, 17)    <= sub_wire237(17);
	sub_wire2(20, 18)    <= sub_wire237(18);
	sub_wire2(20, 19)    <= sub_wire237(19);
	sub_wire2(20, 20)    <= sub_wire237(20);
	sub_wire2(20, 21)    <= sub_wire237(21);
	sub_wire2(20, 22)    <= sub_wire237(22);
	sub_wire2(20, 23)    <= sub_wire237(23);
	sub_wire2(20, 24)    <= sub_wire237(24);
	sub_wire2(20, 25)    <= sub_wire237(25);
	sub_wire2(20, 26)    <= sub_wire237(26);
	sub_wire2(20, 27)    <= sub_wire237(27);
	sub_wire2(20, 28)    <= sub_wire237(28);
	sub_wire2(20, 29)    <= sub_wire237(29);
	sub_wire2(20, 30)    <= sub_wire237(30);
	sub_wire2(20, 31)    <= sub_wire237(31);
	sub_wire2(20, 32)    <= sub_wire237(32);
	sub_wire2(20, 33)    <= sub_wire237(33);
	sub_wire2(20, 34)    <= sub_wire237(34);
	sub_wire2(20, 35)    <= sub_wire237(35);
	sub_wire2(20, 36)    <= sub_wire237(36);
	sub_wire2(20, 37)    <= sub_wire237(37);
	sub_wire2(20, 38)    <= sub_wire237(38);
	sub_wire2(20, 39)    <= sub_wire237(39);
	sub_wire2(19, 0)    <= sub_wire238(0);
	sub_wire2(19, 1)    <= sub_wire238(1);
	sub_wire2(19, 2)    <= sub_wire238(2);
	sub_wire2(19, 3)    <= sub_wire238(3);
	sub_wire2(19, 4)    <= sub_wire238(4);
	sub_wire2(19, 5)    <= sub_wire238(5);
	sub_wire2(19, 6)    <= sub_wire238(6);
	sub_wire2(19, 7)    <= sub_wire238(7);
	sub_wire2(19, 8)    <= sub_wire238(8);
	sub_wire2(19, 9)    <= sub_wire238(9);
	sub_wire2(19, 10)    <= sub_wire238(10);
	sub_wire2(19, 11)    <= sub_wire238(11);
	sub_wire2(19, 12)    <= sub_wire238(12);
	sub_wire2(19, 13)    <= sub_wire238(13);
	sub_wire2(19, 14)    <= sub_wire238(14);
	sub_wire2(19, 15)    <= sub_wire238(15);
	sub_wire2(19, 16)    <= sub_wire238(16);
	sub_wire2(19, 17)    <= sub_wire238(17);
	sub_wire2(19, 18)    <= sub_wire238(18);
	sub_wire2(19, 19)    <= sub_wire238(19);
	sub_wire2(19, 20)    <= sub_wire238(20);
	sub_wire2(19, 21)    <= sub_wire238(21);
	sub_wire2(19, 22)    <= sub_wire238(22);
	sub_wire2(19, 23)    <= sub_wire238(23);
	sub_wire2(19, 24)    <= sub_wire238(24);
	sub_wire2(19, 25)    <= sub_wire238(25);
	sub_wire2(19, 26)    <= sub_wire238(26);
	sub_wire2(19, 27)    <= sub_wire238(27);
	sub_wire2(19, 28)    <= sub_wire238(28);
	sub_wire2(19, 29)    <= sub_wire238(29);
	sub_wire2(19, 30)    <= sub_wire238(30);
	sub_wire2(19, 31)    <= sub_wire238(31);
	sub_wire2(19, 32)    <= sub_wire238(32);
	sub_wire2(19, 33)    <= sub_wire238(33);
	sub_wire2(19, 34)    <= sub_wire238(34);
	sub_wire2(19, 35)    <= sub_wire238(35);
	sub_wire2(19, 36)    <= sub_wire238(36);
	sub_wire2(19, 37)    <= sub_wire238(37);
	sub_wire2(19, 38)    <= sub_wire238(38);
	sub_wire2(19, 39)    <= sub_wire238(39);
	sub_wire2(18, 0)    <= sub_wire239(0);
	sub_wire2(18, 1)    <= sub_wire239(1);
	sub_wire2(18, 2)    <= sub_wire239(2);
	sub_wire2(18, 3)    <= sub_wire239(3);
	sub_wire2(18, 4)    <= sub_wire239(4);
	sub_wire2(18, 5)    <= sub_wire239(5);
	sub_wire2(18, 6)    <= sub_wire239(6);
	sub_wire2(18, 7)    <= sub_wire239(7);
	sub_wire2(18, 8)    <= sub_wire239(8);
	sub_wire2(18, 9)    <= sub_wire239(9);
	sub_wire2(18, 10)    <= sub_wire239(10);
	sub_wire2(18, 11)    <= sub_wire239(11);
	sub_wire2(18, 12)    <= sub_wire239(12);
	sub_wire2(18, 13)    <= sub_wire239(13);
	sub_wire2(18, 14)    <= sub_wire239(14);
	sub_wire2(18, 15)    <= sub_wire239(15);
	sub_wire2(18, 16)    <= sub_wire239(16);
	sub_wire2(18, 17)    <= sub_wire239(17);
	sub_wire2(18, 18)    <= sub_wire239(18);
	sub_wire2(18, 19)    <= sub_wire239(19);
	sub_wire2(18, 20)    <= sub_wire239(20);
	sub_wire2(18, 21)    <= sub_wire239(21);
	sub_wire2(18, 22)    <= sub_wire239(22);
	sub_wire2(18, 23)    <= sub_wire239(23);
	sub_wire2(18, 24)    <= sub_wire239(24);
	sub_wire2(18, 25)    <= sub_wire239(25);
	sub_wire2(18, 26)    <= sub_wire239(26);
	sub_wire2(18, 27)    <= sub_wire239(27);
	sub_wire2(18, 28)    <= sub_wire239(28);
	sub_wire2(18, 29)    <= sub_wire239(29);
	sub_wire2(18, 30)    <= sub_wire239(30);
	sub_wire2(18, 31)    <= sub_wire239(31);
	sub_wire2(18, 32)    <= sub_wire239(32);
	sub_wire2(18, 33)    <= sub_wire239(33);
	sub_wire2(18, 34)    <= sub_wire239(34);
	sub_wire2(18, 35)    <= sub_wire239(35);
	sub_wire2(18, 36)    <= sub_wire239(36);
	sub_wire2(18, 37)    <= sub_wire239(37);
	sub_wire2(18, 38)    <= sub_wire239(38);
	sub_wire2(18, 39)    <= sub_wire239(39);
	sub_wire2(17, 0)    <= sub_wire240(0);
	sub_wire2(17, 1)    <= sub_wire240(1);
	sub_wire2(17, 2)    <= sub_wire240(2);
	sub_wire2(17, 3)    <= sub_wire240(3);
	sub_wire2(17, 4)    <= sub_wire240(4);
	sub_wire2(17, 5)    <= sub_wire240(5);
	sub_wire2(17, 6)    <= sub_wire240(6);
	sub_wire2(17, 7)    <= sub_wire240(7);
	sub_wire2(17, 8)    <= sub_wire240(8);
	sub_wire2(17, 9)    <= sub_wire240(9);
	sub_wire2(17, 10)    <= sub_wire240(10);
	sub_wire2(17, 11)    <= sub_wire240(11);
	sub_wire2(17, 12)    <= sub_wire240(12);
	sub_wire2(17, 13)    <= sub_wire240(13);
	sub_wire2(17, 14)    <= sub_wire240(14);
	sub_wire2(17, 15)    <= sub_wire240(15);
	sub_wire2(17, 16)    <= sub_wire240(16);
	sub_wire2(17, 17)    <= sub_wire240(17);
	sub_wire2(17, 18)    <= sub_wire240(18);
	sub_wire2(17, 19)    <= sub_wire240(19);
	sub_wire2(17, 20)    <= sub_wire240(20);
	sub_wire2(17, 21)    <= sub_wire240(21);
	sub_wire2(17, 22)    <= sub_wire240(22);
	sub_wire2(17, 23)    <= sub_wire240(23);
	sub_wire2(17, 24)    <= sub_wire240(24);
	sub_wire2(17, 25)    <= sub_wire240(25);
	sub_wire2(17, 26)    <= sub_wire240(26);
	sub_wire2(17, 27)    <= sub_wire240(27);
	sub_wire2(17, 28)    <= sub_wire240(28);
	sub_wire2(17, 29)    <= sub_wire240(29);
	sub_wire2(17, 30)    <= sub_wire240(30);
	sub_wire2(17, 31)    <= sub_wire240(31);
	sub_wire2(17, 32)    <= sub_wire240(32);
	sub_wire2(17, 33)    <= sub_wire240(33);
	sub_wire2(17, 34)    <= sub_wire240(34);
	sub_wire2(17, 35)    <= sub_wire240(35);
	sub_wire2(17, 36)    <= sub_wire240(36);
	sub_wire2(17, 37)    <= sub_wire240(37);
	sub_wire2(17, 38)    <= sub_wire240(38);
	sub_wire2(17, 39)    <= sub_wire240(39);
	sub_wire2(16, 0)    <= sub_wire241(0);
	sub_wire2(16, 1)    <= sub_wire241(1);
	sub_wire2(16, 2)    <= sub_wire241(2);
	sub_wire2(16, 3)    <= sub_wire241(3);
	sub_wire2(16, 4)    <= sub_wire241(4);
	sub_wire2(16, 5)    <= sub_wire241(5);
	sub_wire2(16, 6)    <= sub_wire241(6);
	sub_wire2(16, 7)    <= sub_wire241(7);
	sub_wire2(16, 8)    <= sub_wire241(8);
	sub_wire2(16, 9)    <= sub_wire241(9);
	sub_wire2(16, 10)    <= sub_wire241(10);
	sub_wire2(16, 11)    <= sub_wire241(11);
	sub_wire2(16, 12)    <= sub_wire241(12);
	sub_wire2(16, 13)    <= sub_wire241(13);
	sub_wire2(16, 14)    <= sub_wire241(14);
	sub_wire2(16, 15)    <= sub_wire241(15);
	sub_wire2(16, 16)    <= sub_wire241(16);
	sub_wire2(16, 17)    <= sub_wire241(17);
	sub_wire2(16, 18)    <= sub_wire241(18);
	sub_wire2(16, 19)    <= sub_wire241(19);
	sub_wire2(16, 20)    <= sub_wire241(20);
	sub_wire2(16, 21)    <= sub_wire241(21);
	sub_wire2(16, 22)    <= sub_wire241(22);
	sub_wire2(16, 23)    <= sub_wire241(23);
	sub_wire2(16, 24)    <= sub_wire241(24);
	sub_wire2(16, 25)    <= sub_wire241(25);
	sub_wire2(16, 26)    <= sub_wire241(26);
	sub_wire2(16, 27)    <= sub_wire241(27);
	sub_wire2(16, 28)    <= sub_wire241(28);
	sub_wire2(16, 29)    <= sub_wire241(29);
	sub_wire2(16, 30)    <= sub_wire241(30);
	sub_wire2(16, 31)    <= sub_wire241(31);
	sub_wire2(16, 32)    <= sub_wire241(32);
	sub_wire2(16, 33)    <= sub_wire241(33);
	sub_wire2(16, 34)    <= sub_wire241(34);
	sub_wire2(16, 35)    <= sub_wire241(35);
	sub_wire2(16, 36)    <= sub_wire241(36);
	sub_wire2(16, 37)    <= sub_wire241(37);
	sub_wire2(16, 38)    <= sub_wire241(38);
	sub_wire2(16, 39)    <= sub_wire241(39);
	sub_wire2(15, 0)    <= sub_wire242(0);
	sub_wire2(15, 1)    <= sub_wire242(1);
	sub_wire2(15, 2)    <= sub_wire242(2);
	sub_wire2(15, 3)    <= sub_wire242(3);
	sub_wire2(15, 4)    <= sub_wire242(4);
	sub_wire2(15, 5)    <= sub_wire242(5);
	sub_wire2(15, 6)    <= sub_wire242(6);
	sub_wire2(15, 7)    <= sub_wire242(7);
	sub_wire2(15, 8)    <= sub_wire242(8);
	sub_wire2(15, 9)    <= sub_wire242(9);
	sub_wire2(15, 10)    <= sub_wire242(10);
	sub_wire2(15, 11)    <= sub_wire242(11);
	sub_wire2(15, 12)    <= sub_wire242(12);
	sub_wire2(15, 13)    <= sub_wire242(13);
	sub_wire2(15, 14)    <= sub_wire242(14);
	sub_wire2(15, 15)    <= sub_wire242(15);
	sub_wire2(15, 16)    <= sub_wire242(16);
	sub_wire2(15, 17)    <= sub_wire242(17);
	sub_wire2(15, 18)    <= sub_wire242(18);
	sub_wire2(15, 19)    <= sub_wire242(19);
	sub_wire2(15, 20)    <= sub_wire242(20);
	sub_wire2(15, 21)    <= sub_wire242(21);
	sub_wire2(15, 22)    <= sub_wire242(22);
	sub_wire2(15, 23)    <= sub_wire242(23);
	sub_wire2(15, 24)    <= sub_wire242(24);
	sub_wire2(15, 25)    <= sub_wire242(25);
	sub_wire2(15, 26)    <= sub_wire242(26);
	sub_wire2(15, 27)    <= sub_wire242(27);
	sub_wire2(15, 28)    <= sub_wire242(28);
	sub_wire2(15, 29)    <= sub_wire242(29);
	sub_wire2(15, 30)    <= sub_wire242(30);
	sub_wire2(15, 31)    <= sub_wire242(31);
	sub_wire2(15, 32)    <= sub_wire242(32);
	sub_wire2(15, 33)    <= sub_wire242(33);
	sub_wire2(15, 34)    <= sub_wire242(34);
	sub_wire2(15, 35)    <= sub_wire242(35);
	sub_wire2(15, 36)    <= sub_wire242(36);
	sub_wire2(15, 37)    <= sub_wire242(37);
	sub_wire2(15, 38)    <= sub_wire242(38);
	sub_wire2(15, 39)    <= sub_wire242(39);
	sub_wire2(14, 0)    <= sub_wire243(0);
	sub_wire2(14, 1)    <= sub_wire243(1);
	sub_wire2(14, 2)    <= sub_wire243(2);
	sub_wire2(14, 3)    <= sub_wire243(3);
	sub_wire2(14, 4)    <= sub_wire243(4);
	sub_wire2(14, 5)    <= sub_wire243(5);
	sub_wire2(14, 6)    <= sub_wire243(6);
	sub_wire2(14, 7)    <= sub_wire243(7);
	sub_wire2(14, 8)    <= sub_wire243(8);
	sub_wire2(14, 9)    <= sub_wire243(9);
	sub_wire2(14, 10)    <= sub_wire243(10);
	sub_wire2(14, 11)    <= sub_wire243(11);
	sub_wire2(14, 12)    <= sub_wire243(12);
	sub_wire2(14, 13)    <= sub_wire243(13);
	sub_wire2(14, 14)    <= sub_wire243(14);
	sub_wire2(14, 15)    <= sub_wire243(15);
	sub_wire2(14, 16)    <= sub_wire243(16);
	sub_wire2(14, 17)    <= sub_wire243(17);
	sub_wire2(14, 18)    <= sub_wire243(18);
	sub_wire2(14, 19)    <= sub_wire243(19);
	sub_wire2(14, 20)    <= sub_wire243(20);
	sub_wire2(14, 21)    <= sub_wire243(21);
	sub_wire2(14, 22)    <= sub_wire243(22);
	sub_wire2(14, 23)    <= sub_wire243(23);
	sub_wire2(14, 24)    <= sub_wire243(24);
	sub_wire2(14, 25)    <= sub_wire243(25);
	sub_wire2(14, 26)    <= sub_wire243(26);
	sub_wire2(14, 27)    <= sub_wire243(27);
	sub_wire2(14, 28)    <= sub_wire243(28);
	sub_wire2(14, 29)    <= sub_wire243(29);
	sub_wire2(14, 30)    <= sub_wire243(30);
	sub_wire2(14, 31)    <= sub_wire243(31);
	sub_wire2(14, 32)    <= sub_wire243(32);
	sub_wire2(14, 33)    <= sub_wire243(33);
	sub_wire2(14, 34)    <= sub_wire243(34);
	sub_wire2(14, 35)    <= sub_wire243(35);
	sub_wire2(14, 36)    <= sub_wire243(36);
	sub_wire2(14, 37)    <= sub_wire243(37);
	sub_wire2(14, 38)    <= sub_wire243(38);
	sub_wire2(14, 39)    <= sub_wire243(39);
	sub_wire2(13, 0)    <= sub_wire244(0);
	sub_wire2(13, 1)    <= sub_wire244(1);
	sub_wire2(13, 2)    <= sub_wire244(2);
	sub_wire2(13, 3)    <= sub_wire244(3);
	sub_wire2(13, 4)    <= sub_wire244(4);
	sub_wire2(13, 5)    <= sub_wire244(5);
	sub_wire2(13, 6)    <= sub_wire244(6);
	sub_wire2(13, 7)    <= sub_wire244(7);
	sub_wire2(13, 8)    <= sub_wire244(8);
	sub_wire2(13, 9)    <= sub_wire244(9);
	sub_wire2(13, 10)    <= sub_wire244(10);
	sub_wire2(13, 11)    <= sub_wire244(11);
	sub_wire2(13, 12)    <= sub_wire244(12);
	sub_wire2(13, 13)    <= sub_wire244(13);
	sub_wire2(13, 14)    <= sub_wire244(14);
	sub_wire2(13, 15)    <= sub_wire244(15);
	sub_wire2(13, 16)    <= sub_wire244(16);
	sub_wire2(13, 17)    <= sub_wire244(17);
	sub_wire2(13, 18)    <= sub_wire244(18);
	sub_wire2(13, 19)    <= sub_wire244(19);
	sub_wire2(13, 20)    <= sub_wire244(20);
	sub_wire2(13, 21)    <= sub_wire244(21);
	sub_wire2(13, 22)    <= sub_wire244(22);
	sub_wire2(13, 23)    <= sub_wire244(23);
	sub_wire2(13, 24)    <= sub_wire244(24);
	sub_wire2(13, 25)    <= sub_wire244(25);
	sub_wire2(13, 26)    <= sub_wire244(26);
	sub_wire2(13, 27)    <= sub_wire244(27);
	sub_wire2(13, 28)    <= sub_wire244(28);
	sub_wire2(13, 29)    <= sub_wire244(29);
	sub_wire2(13, 30)    <= sub_wire244(30);
	sub_wire2(13, 31)    <= sub_wire244(31);
	sub_wire2(13, 32)    <= sub_wire244(32);
	sub_wire2(13, 33)    <= sub_wire244(33);
	sub_wire2(13, 34)    <= sub_wire244(34);
	sub_wire2(13, 35)    <= sub_wire244(35);
	sub_wire2(13, 36)    <= sub_wire244(36);
	sub_wire2(13, 37)    <= sub_wire244(37);
	sub_wire2(13, 38)    <= sub_wire244(38);
	sub_wire2(13, 39)    <= sub_wire244(39);
	sub_wire2(12, 0)    <= sub_wire245(0);
	sub_wire2(12, 1)    <= sub_wire245(1);
	sub_wire2(12, 2)    <= sub_wire245(2);
	sub_wire2(12, 3)    <= sub_wire245(3);
	sub_wire2(12, 4)    <= sub_wire245(4);
	sub_wire2(12, 5)    <= sub_wire245(5);
	sub_wire2(12, 6)    <= sub_wire245(6);
	sub_wire2(12, 7)    <= sub_wire245(7);
	sub_wire2(12, 8)    <= sub_wire245(8);
	sub_wire2(12, 9)    <= sub_wire245(9);
	sub_wire2(12, 10)    <= sub_wire245(10);
	sub_wire2(12, 11)    <= sub_wire245(11);
	sub_wire2(12, 12)    <= sub_wire245(12);
	sub_wire2(12, 13)    <= sub_wire245(13);
	sub_wire2(12, 14)    <= sub_wire245(14);
	sub_wire2(12, 15)    <= sub_wire245(15);
	sub_wire2(12, 16)    <= sub_wire245(16);
	sub_wire2(12, 17)    <= sub_wire245(17);
	sub_wire2(12, 18)    <= sub_wire245(18);
	sub_wire2(12, 19)    <= sub_wire245(19);
	sub_wire2(12, 20)    <= sub_wire245(20);
	sub_wire2(12, 21)    <= sub_wire245(21);
	sub_wire2(12, 22)    <= sub_wire245(22);
	sub_wire2(12, 23)    <= sub_wire245(23);
	sub_wire2(12, 24)    <= sub_wire245(24);
	sub_wire2(12, 25)    <= sub_wire245(25);
	sub_wire2(12, 26)    <= sub_wire245(26);
	sub_wire2(12, 27)    <= sub_wire245(27);
	sub_wire2(12, 28)    <= sub_wire245(28);
	sub_wire2(12, 29)    <= sub_wire245(29);
	sub_wire2(12, 30)    <= sub_wire245(30);
	sub_wire2(12, 31)    <= sub_wire245(31);
	sub_wire2(12, 32)    <= sub_wire245(32);
	sub_wire2(12, 33)    <= sub_wire245(33);
	sub_wire2(12, 34)    <= sub_wire245(34);
	sub_wire2(12, 35)    <= sub_wire245(35);
	sub_wire2(12, 36)    <= sub_wire245(36);
	sub_wire2(12, 37)    <= sub_wire245(37);
	sub_wire2(12, 38)    <= sub_wire245(38);
	sub_wire2(12, 39)    <= sub_wire245(39);
	sub_wire2(11, 0)    <= sub_wire246(0);
	sub_wire2(11, 1)    <= sub_wire246(1);
	sub_wire2(11, 2)    <= sub_wire246(2);
	sub_wire2(11, 3)    <= sub_wire246(3);
	sub_wire2(11, 4)    <= sub_wire246(4);
	sub_wire2(11, 5)    <= sub_wire246(5);
	sub_wire2(11, 6)    <= sub_wire246(6);
	sub_wire2(11, 7)    <= sub_wire246(7);
	sub_wire2(11, 8)    <= sub_wire246(8);
	sub_wire2(11, 9)    <= sub_wire246(9);
	sub_wire2(11, 10)    <= sub_wire246(10);
	sub_wire2(11, 11)    <= sub_wire246(11);
	sub_wire2(11, 12)    <= sub_wire246(12);
	sub_wire2(11, 13)    <= sub_wire246(13);
	sub_wire2(11, 14)    <= sub_wire246(14);
	sub_wire2(11, 15)    <= sub_wire246(15);
	sub_wire2(11, 16)    <= sub_wire246(16);
	sub_wire2(11, 17)    <= sub_wire246(17);
	sub_wire2(11, 18)    <= sub_wire246(18);
	sub_wire2(11, 19)    <= sub_wire246(19);
	sub_wire2(11, 20)    <= sub_wire246(20);
	sub_wire2(11, 21)    <= sub_wire246(21);
	sub_wire2(11, 22)    <= sub_wire246(22);
	sub_wire2(11, 23)    <= sub_wire246(23);
	sub_wire2(11, 24)    <= sub_wire246(24);
	sub_wire2(11, 25)    <= sub_wire246(25);
	sub_wire2(11, 26)    <= sub_wire246(26);
	sub_wire2(11, 27)    <= sub_wire246(27);
	sub_wire2(11, 28)    <= sub_wire246(28);
	sub_wire2(11, 29)    <= sub_wire246(29);
	sub_wire2(11, 30)    <= sub_wire246(30);
	sub_wire2(11, 31)    <= sub_wire246(31);
	sub_wire2(11, 32)    <= sub_wire246(32);
	sub_wire2(11, 33)    <= sub_wire246(33);
	sub_wire2(11, 34)    <= sub_wire246(34);
	sub_wire2(11, 35)    <= sub_wire246(35);
	sub_wire2(11, 36)    <= sub_wire246(36);
	sub_wire2(11, 37)    <= sub_wire246(37);
	sub_wire2(11, 38)    <= sub_wire246(38);
	sub_wire2(11, 39)    <= sub_wire246(39);
	sub_wire2(10, 0)    <= sub_wire247(0);
	sub_wire2(10, 1)    <= sub_wire247(1);
	sub_wire2(10, 2)    <= sub_wire247(2);
	sub_wire2(10, 3)    <= sub_wire247(3);
	sub_wire2(10, 4)    <= sub_wire247(4);
	sub_wire2(10, 5)    <= sub_wire247(5);
	sub_wire2(10, 6)    <= sub_wire247(6);
	sub_wire2(10, 7)    <= sub_wire247(7);
	sub_wire2(10, 8)    <= sub_wire247(8);
	sub_wire2(10, 9)    <= sub_wire247(9);
	sub_wire2(10, 10)    <= sub_wire247(10);
	sub_wire2(10, 11)    <= sub_wire247(11);
	sub_wire2(10, 12)    <= sub_wire247(12);
	sub_wire2(10, 13)    <= sub_wire247(13);
	sub_wire2(10, 14)    <= sub_wire247(14);
	sub_wire2(10, 15)    <= sub_wire247(15);
	sub_wire2(10, 16)    <= sub_wire247(16);
	sub_wire2(10, 17)    <= sub_wire247(17);
	sub_wire2(10, 18)    <= sub_wire247(18);
	sub_wire2(10, 19)    <= sub_wire247(19);
	sub_wire2(10, 20)    <= sub_wire247(20);
	sub_wire2(10, 21)    <= sub_wire247(21);
	sub_wire2(10, 22)    <= sub_wire247(22);
	sub_wire2(10, 23)    <= sub_wire247(23);
	sub_wire2(10, 24)    <= sub_wire247(24);
	sub_wire2(10, 25)    <= sub_wire247(25);
	sub_wire2(10, 26)    <= sub_wire247(26);
	sub_wire2(10, 27)    <= sub_wire247(27);
	sub_wire2(10, 28)    <= sub_wire247(28);
	sub_wire2(10, 29)    <= sub_wire247(29);
	sub_wire2(10, 30)    <= sub_wire247(30);
	sub_wire2(10, 31)    <= sub_wire247(31);
	sub_wire2(10, 32)    <= sub_wire247(32);
	sub_wire2(10, 33)    <= sub_wire247(33);
	sub_wire2(10, 34)    <= sub_wire247(34);
	sub_wire2(10, 35)    <= sub_wire247(35);
	sub_wire2(10, 36)    <= sub_wire247(36);
	sub_wire2(10, 37)    <= sub_wire247(37);
	sub_wire2(10, 38)    <= sub_wire247(38);
	sub_wire2(10, 39)    <= sub_wire247(39);
	sub_wire2(9, 0)    <= sub_wire248(0);
	sub_wire2(9, 1)    <= sub_wire248(1);
	sub_wire2(9, 2)    <= sub_wire248(2);
	sub_wire2(9, 3)    <= sub_wire248(3);
	sub_wire2(9, 4)    <= sub_wire248(4);
	sub_wire2(9, 5)    <= sub_wire248(5);
	sub_wire2(9, 6)    <= sub_wire248(6);
	sub_wire2(9, 7)    <= sub_wire248(7);
	sub_wire2(9, 8)    <= sub_wire248(8);
	sub_wire2(9, 9)    <= sub_wire248(9);
	sub_wire2(9, 10)    <= sub_wire248(10);
	sub_wire2(9, 11)    <= sub_wire248(11);
	sub_wire2(9, 12)    <= sub_wire248(12);
	sub_wire2(9, 13)    <= sub_wire248(13);
	sub_wire2(9, 14)    <= sub_wire248(14);
	sub_wire2(9, 15)    <= sub_wire248(15);
	sub_wire2(9, 16)    <= sub_wire248(16);
	sub_wire2(9, 17)    <= sub_wire248(17);
	sub_wire2(9, 18)    <= sub_wire248(18);
	sub_wire2(9, 19)    <= sub_wire248(19);
	sub_wire2(9, 20)    <= sub_wire248(20);
	sub_wire2(9, 21)    <= sub_wire248(21);
	sub_wire2(9, 22)    <= sub_wire248(22);
	sub_wire2(9, 23)    <= sub_wire248(23);
	sub_wire2(9, 24)    <= sub_wire248(24);
	sub_wire2(9, 25)    <= sub_wire248(25);
	sub_wire2(9, 26)    <= sub_wire248(26);
	sub_wire2(9, 27)    <= sub_wire248(27);
	sub_wire2(9, 28)    <= sub_wire248(28);
	sub_wire2(9, 29)    <= sub_wire248(29);
	sub_wire2(9, 30)    <= sub_wire248(30);
	sub_wire2(9, 31)    <= sub_wire248(31);
	sub_wire2(9, 32)    <= sub_wire248(32);
	sub_wire2(9, 33)    <= sub_wire248(33);
	sub_wire2(9, 34)    <= sub_wire248(34);
	sub_wire2(9, 35)    <= sub_wire248(35);
	sub_wire2(9, 36)    <= sub_wire248(36);
	sub_wire2(9, 37)    <= sub_wire248(37);
	sub_wire2(9, 38)    <= sub_wire248(38);
	sub_wire2(9, 39)    <= sub_wire248(39);
	sub_wire2(8, 0)    <= sub_wire249(0);
	sub_wire2(8, 1)    <= sub_wire249(1);
	sub_wire2(8, 2)    <= sub_wire249(2);
	sub_wire2(8, 3)    <= sub_wire249(3);
	sub_wire2(8, 4)    <= sub_wire249(4);
	sub_wire2(8, 5)    <= sub_wire249(5);
	sub_wire2(8, 6)    <= sub_wire249(6);
	sub_wire2(8, 7)    <= sub_wire249(7);
	sub_wire2(8, 8)    <= sub_wire249(8);
	sub_wire2(8, 9)    <= sub_wire249(9);
	sub_wire2(8, 10)    <= sub_wire249(10);
	sub_wire2(8, 11)    <= sub_wire249(11);
	sub_wire2(8, 12)    <= sub_wire249(12);
	sub_wire2(8, 13)    <= sub_wire249(13);
	sub_wire2(8, 14)    <= sub_wire249(14);
	sub_wire2(8, 15)    <= sub_wire249(15);
	sub_wire2(8, 16)    <= sub_wire249(16);
	sub_wire2(8, 17)    <= sub_wire249(17);
	sub_wire2(8, 18)    <= sub_wire249(18);
	sub_wire2(8, 19)    <= sub_wire249(19);
	sub_wire2(8, 20)    <= sub_wire249(20);
	sub_wire2(8, 21)    <= sub_wire249(21);
	sub_wire2(8, 22)    <= sub_wire249(22);
	sub_wire2(8, 23)    <= sub_wire249(23);
	sub_wire2(8, 24)    <= sub_wire249(24);
	sub_wire2(8, 25)    <= sub_wire249(25);
	sub_wire2(8, 26)    <= sub_wire249(26);
	sub_wire2(8, 27)    <= sub_wire249(27);
	sub_wire2(8, 28)    <= sub_wire249(28);
	sub_wire2(8, 29)    <= sub_wire249(29);
	sub_wire2(8, 30)    <= sub_wire249(30);
	sub_wire2(8, 31)    <= sub_wire249(31);
	sub_wire2(8, 32)    <= sub_wire249(32);
	sub_wire2(8, 33)    <= sub_wire249(33);
	sub_wire2(8, 34)    <= sub_wire249(34);
	sub_wire2(8, 35)    <= sub_wire249(35);
	sub_wire2(8, 36)    <= sub_wire249(36);
	sub_wire2(8, 37)    <= sub_wire249(37);
	sub_wire2(8, 38)    <= sub_wire249(38);
	sub_wire2(8, 39)    <= sub_wire249(39);
	sub_wire2(7, 0)    <= sub_wire250(0);
	sub_wire2(7, 1)    <= sub_wire250(1);
	sub_wire2(7, 2)    <= sub_wire250(2);
	sub_wire2(7, 3)    <= sub_wire250(3);
	sub_wire2(7, 4)    <= sub_wire250(4);
	sub_wire2(7, 5)    <= sub_wire250(5);
	sub_wire2(7, 6)    <= sub_wire250(6);
	sub_wire2(7, 7)    <= sub_wire250(7);
	sub_wire2(7, 8)    <= sub_wire250(8);
	sub_wire2(7, 9)    <= sub_wire250(9);
	sub_wire2(7, 10)    <= sub_wire250(10);
	sub_wire2(7, 11)    <= sub_wire250(11);
	sub_wire2(7, 12)    <= sub_wire250(12);
	sub_wire2(7, 13)    <= sub_wire250(13);
	sub_wire2(7, 14)    <= sub_wire250(14);
	sub_wire2(7, 15)    <= sub_wire250(15);
	sub_wire2(7, 16)    <= sub_wire250(16);
	sub_wire2(7, 17)    <= sub_wire250(17);
	sub_wire2(7, 18)    <= sub_wire250(18);
	sub_wire2(7, 19)    <= sub_wire250(19);
	sub_wire2(7, 20)    <= sub_wire250(20);
	sub_wire2(7, 21)    <= sub_wire250(21);
	sub_wire2(7, 22)    <= sub_wire250(22);
	sub_wire2(7, 23)    <= sub_wire250(23);
	sub_wire2(7, 24)    <= sub_wire250(24);
	sub_wire2(7, 25)    <= sub_wire250(25);
	sub_wire2(7, 26)    <= sub_wire250(26);
	sub_wire2(7, 27)    <= sub_wire250(27);
	sub_wire2(7, 28)    <= sub_wire250(28);
	sub_wire2(7, 29)    <= sub_wire250(29);
	sub_wire2(7, 30)    <= sub_wire250(30);
	sub_wire2(7, 31)    <= sub_wire250(31);
	sub_wire2(7, 32)    <= sub_wire250(32);
	sub_wire2(7, 33)    <= sub_wire250(33);
	sub_wire2(7, 34)    <= sub_wire250(34);
	sub_wire2(7, 35)    <= sub_wire250(35);
	sub_wire2(7, 36)    <= sub_wire250(36);
	sub_wire2(7, 37)    <= sub_wire250(37);
	sub_wire2(7, 38)    <= sub_wire250(38);
	sub_wire2(7, 39)    <= sub_wire250(39);
	sub_wire2(6, 0)    <= sub_wire251(0);
	sub_wire2(6, 1)    <= sub_wire251(1);
	sub_wire2(6, 2)    <= sub_wire251(2);
	sub_wire2(6, 3)    <= sub_wire251(3);
	sub_wire2(6, 4)    <= sub_wire251(4);
	sub_wire2(6, 5)    <= sub_wire251(5);
	sub_wire2(6, 6)    <= sub_wire251(6);
	sub_wire2(6, 7)    <= sub_wire251(7);
	sub_wire2(6, 8)    <= sub_wire251(8);
	sub_wire2(6, 9)    <= sub_wire251(9);
	sub_wire2(6, 10)    <= sub_wire251(10);
	sub_wire2(6, 11)    <= sub_wire251(11);
	sub_wire2(6, 12)    <= sub_wire251(12);
	sub_wire2(6, 13)    <= sub_wire251(13);
	sub_wire2(6, 14)    <= sub_wire251(14);
	sub_wire2(6, 15)    <= sub_wire251(15);
	sub_wire2(6, 16)    <= sub_wire251(16);
	sub_wire2(6, 17)    <= sub_wire251(17);
	sub_wire2(6, 18)    <= sub_wire251(18);
	sub_wire2(6, 19)    <= sub_wire251(19);
	sub_wire2(6, 20)    <= sub_wire251(20);
	sub_wire2(6, 21)    <= sub_wire251(21);
	sub_wire2(6, 22)    <= sub_wire251(22);
	sub_wire2(6, 23)    <= sub_wire251(23);
	sub_wire2(6, 24)    <= sub_wire251(24);
	sub_wire2(6, 25)    <= sub_wire251(25);
	sub_wire2(6, 26)    <= sub_wire251(26);
	sub_wire2(6, 27)    <= sub_wire251(27);
	sub_wire2(6, 28)    <= sub_wire251(28);
	sub_wire2(6, 29)    <= sub_wire251(29);
	sub_wire2(6, 30)    <= sub_wire251(30);
	sub_wire2(6, 31)    <= sub_wire251(31);
	sub_wire2(6, 32)    <= sub_wire251(32);
	sub_wire2(6, 33)    <= sub_wire251(33);
	sub_wire2(6, 34)    <= sub_wire251(34);
	sub_wire2(6, 35)    <= sub_wire251(35);
	sub_wire2(6, 36)    <= sub_wire251(36);
	sub_wire2(6, 37)    <= sub_wire251(37);
	sub_wire2(6, 38)    <= sub_wire251(38);
	sub_wire2(6, 39)    <= sub_wire251(39);
	sub_wire2(5, 0)    <= sub_wire252(0);
	sub_wire2(5, 1)    <= sub_wire252(1);
	sub_wire2(5, 2)    <= sub_wire252(2);
	sub_wire2(5, 3)    <= sub_wire252(3);
	sub_wire2(5, 4)    <= sub_wire252(4);
	sub_wire2(5, 5)    <= sub_wire252(5);
	sub_wire2(5, 6)    <= sub_wire252(6);
	sub_wire2(5, 7)    <= sub_wire252(7);
	sub_wire2(5, 8)    <= sub_wire252(8);
	sub_wire2(5, 9)    <= sub_wire252(9);
	sub_wire2(5, 10)    <= sub_wire252(10);
	sub_wire2(5, 11)    <= sub_wire252(11);
	sub_wire2(5, 12)    <= sub_wire252(12);
	sub_wire2(5, 13)    <= sub_wire252(13);
	sub_wire2(5, 14)    <= sub_wire252(14);
	sub_wire2(5, 15)    <= sub_wire252(15);
	sub_wire2(5, 16)    <= sub_wire252(16);
	sub_wire2(5, 17)    <= sub_wire252(17);
	sub_wire2(5, 18)    <= sub_wire252(18);
	sub_wire2(5, 19)    <= sub_wire252(19);
	sub_wire2(5, 20)    <= sub_wire252(20);
	sub_wire2(5, 21)    <= sub_wire252(21);
	sub_wire2(5, 22)    <= sub_wire252(22);
	sub_wire2(5, 23)    <= sub_wire252(23);
	sub_wire2(5, 24)    <= sub_wire252(24);
	sub_wire2(5, 25)    <= sub_wire252(25);
	sub_wire2(5, 26)    <= sub_wire252(26);
	sub_wire2(5, 27)    <= sub_wire252(27);
	sub_wire2(5, 28)    <= sub_wire252(28);
	sub_wire2(5, 29)    <= sub_wire252(29);
	sub_wire2(5, 30)    <= sub_wire252(30);
	sub_wire2(5, 31)    <= sub_wire252(31);
	sub_wire2(5, 32)    <= sub_wire252(32);
	sub_wire2(5, 33)    <= sub_wire252(33);
	sub_wire2(5, 34)    <= sub_wire252(34);
	sub_wire2(5, 35)    <= sub_wire252(35);
	sub_wire2(5, 36)    <= sub_wire252(36);
	sub_wire2(5, 37)    <= sub_wire252(37);
	sub_wire2(5, 38)    <= sub_wire252(38);
	sub_wire2(5, 39)    <= sub_wire252(39);
	sub_wire2(4, 0)    <= sub_wire253(0);
	sub_wire2(4, 1)    <= sub_wire253(1);
	sub_wire2(4, 2)    <= sub_wire253(2);
	sub_wire2(4, 3)    <= sub_wire253(3);
	sub_wire2(4, 4)    <= sub_wire253(4);
	sub_wire2(4, 5)    <= sub_wire253(5);
	sub_wire2(4, 6)    <= sub_wire253(6);
	sub_wire2(4, 7)    <= sub_wire253(7);
	sub_wire2(4, 8)    <= sub_wire253(8);
	sub_wire2(4, 9)    <= sub_wire253(9);
	sub_wire2(4, 10)    <= sub_wire253(10);
	sub_wire2(4, 11)    <= sub_wire253(11);
	sub_wire2(4, 12)    <= sub_wire253(12);
	sub_wire2(4, 13)    <= sub_wire253(13);
	sub_wire2(4, 14)    <= sub_wire253(14);
	sub_wire2(4, 15)    <= sub_wire253(15);
	sub_wire2(4, 16)    <= sub_wire253(16);
	sub_wire2(4, 17)    <= sub_wire253(17);
	sub_wire2(4, 18)    <= sub_wire253(18);
	sub_wire2(4, 19)    <= sub_wire253(19);
	sub_wire2(4, 20)    <= sub_wire253(20);
	sub_wire2(4, 21)    <= sub_wire253(21);
	sub_wire2(4, 22)    <= sub_wire253(22);
	sub_wire2(4, 23)    <= sub_wire253(23);
	sub_wire2(4, 24)    <= sub_wire253(24);
	sub_wire2(4, 25)    <= sub_wire253(25);
	sub_wire2(4, 26)    <= sub_wire253(26);
	sub_wire2(4, 27)    <= sub_wire253(27);
	sub_wire2(4, 28)    <= sub_wire253(28);
	sub_wire2(4, 29)    <= sub_wire253(29);
	sub_wire2(4, 30)    <= sub_wire253(30);
	sub_wire2(4, 31)    <= sub_wire253(31);
	sub_wire2(4, 32)    <= sub_wire253(32);
	sub_wire2(4, 33)    <= sub_wire253(33);
	sub_wire2(4, 34)    <= sub_wire253(34);
	sub_wire2(4, 35)    <= sub_wire253(35);
	sub_wire2(4, 36)    <= sub_wire253(36);
	sub_wire2(4, 37)    <= sub_wire253(37);
	sub_wire2(4, 38)    <= sub_wire253(38);
	sub_wire2(4, 39)    <= sub_wire253(39);
	sub_wire2(3, 0)    <= sub_wire254(0);
	sub_wire2(3, 1)    <= sub_wire254(1);
	sub_wire2(3, 2)    <= sub_wire254(2);
	sub_wire2(3, 3)    <= sub_wire254(3);
	sub_wire2(3, 4)    <= sub_wire254(4);
	sub_wire2(3, 5)    <= sub_wire254(5);
	sub_wire2(3, 6)    <= sub_wire254(6);
	sub_wire2(3, 7)    <= sub_wire254(7);
	sub_wire2(3, 8)    <= sub_wire254(8);
	sub_wire2(3, 9)    <= sub_wire254(9);
	sub_wire2(3, 10)    <= sub_wire254(10);
	sub_wire2(3, 11)    <= sub_wire254(11);
	sub_wire2(3, 12)    <= sub_wire254(12);
	sub_wire2(3, 13)    <= sub_wire254(13);
	sub_wire2(3, 14)    <= sub_wire254(14);
	sub_wire2(3, 15)    <= sub_wire254(15);
	sub_wire2(3, 16)    <= sub_wire254(16);
	sub_wire2(3, 17)    <= sub_wire254(17);
	sub_wire2(3, 18)    <= sub_wire254(18);
	sub_wire2(3, 19)    <= sub_wire254(19);
	sub_wire2(3, 20)    <= sub_wire254(20);
	sub_wire2(3, 21)    <= sub_wire254(21);
	sub_wire2(3, 22)    <= sub_wire254(22);
	sub_wire2(3, 23)    <= sub_wire254(23);
	sub_wire2(3, 24)    <= sub_wire254(24);
	sub_wire2(3, 25)    <= sub_wire254(25);
	sub_wire2(3, 26)    <= sub_wire254(26);
	sub_wire2(3, 27)    <= sub_wire254(27);
	sub_wire2(3, 28)    <= sub_wire254(28);
	sub_wire2(3, 29)    <= sub_wire254(29);
	sub_wire2(3, 30)    <= sub_wire254(30);
	sub_wire2(3, 31)    <= sub_wire254(31);
	sub_wire2(3, 32)    <= sub_wire254(32);
	sub_wire2(3, 33)    <= sub_wire254(33);
	sub_wire2(3, 34)    <= sub_wire254(34);
	sub_wire2(3, 35)    <= sub_wire254(35);
	sub_wire2(3, 36)    <= sub_wire254(36);
	sub_wire2(3, 37)    <= sub_wire254(37);
	sub_wire2(3, 38)    <= sub_wire254(38);
	sub_wire2(3, 39)    <= sub_wire254(39);
	sub_wire2(2, 0)    <= sub_wire255(0);
	sub_wire2(2, 1)    <= sub_wire255(1);
	sub_wire2(2, 2)    <= sub_wire255(2);
	sub_wire2(2, 3)    <= sub_wire255(3);
	sub_wire2(2, 4)    <= sub_wire255(4);
	sub_wire2(2, 5)    <= sub_wire255(5);
	sub_wire2(2, 6)    <= sub_wire255(6);
	sub_wire2(2, 7)    <= sub_wire255(7);
	sub_wire2(2, 8)    <= sub_wire255(8);
	sub_wire2(2, 9)    <= sub_wire255(9);
	sub_wire2(2, 10)    <= sub_wire255(10);
	sub_wire2(2, 11)    <= sub_wire255(11);
	sub_wire2(2, 12)    <= sub_wire255(12);
	sub_wire2(2, 13)    <= sub_wire255(13);
	sub_wire2(2, 14)    <= sub_wire255(14);
	sub_wire2(2, 15)    <= sub_wire255(15);
	sub_wire2(2, 16)    <= sub_wire255(16);
	sub_wire2(2, 17)    <= sub_wire255(17);
	sub_wire2(2, 18)    <= sub_wire255(18);
	sub_wire2(2, 19)    <= sub_wire255(19);
	sub_wire2(2, 20)    <= sub_wire255(20);
	sub_wire2(2, 21)    <= sub_wire255(21);
	sub_wire2(2, 22)    <= sub_wire255(22);
	sub_wire2(2, 23)    <= sub_wire255(23);
	sub_wire2(2, 24)    <= sub_wire255(24);
	sub_wire2(2, 25)    <= sub_wire255(25);
	sub_wire2(2, 26)    <= sub_wire255(26);
	sub_wire2(2, 27)    <= sub_wire255(27);
	sub_wire2(2, 28)    <= sub_wire255(28);
	sub_wire2(2, 29)    <= sub_wire255(29);
	sub_wire2(2, 30)    <= sub_wire255(30);
	sub_wire2(2, 31)    <= sub_wire255(31);
	sub_wire2(2, 32)    <= sub_wire255(32);
	sub_wire2(2, 33)    <= sub_wire255(33);
	sub_wire2(2, 34)    <= sub_wire255(34);
	sub_wire2(2, 35)    <= sub_wire255(35);
	sub_wire2(2, 36)    <= sub_wire255(36);
	sub_wire2(2, 37)    <= sub_wire255(37);
	sub_wire2(2, 38)    <= sub_wire255(38);
	sub_wire2(2, 39)    <= sub_wire255(39);
	sub_wire2(1, 0)    <= sub_wire256(0);
	sub_wire2(1, 1)    <= sub_wire256(1);
	sub_wire2(1, 2)    <= sub_wire256(2);
	sub_wire2(1, 3)    <= sub_wire256(3);
	sub_wire2(1, 4)    <= sub_wire256(4);
	sub_wire2(1, 5)    <= sub_wire256(5);
	sub_wire2(1, 6)    <= sub_wire256(6);
	sub_wire2(1, 7)    <= sub_wire256(7);
	sub_wire2(1, 8)    <= sub_wire256(8);
	sub_wire2(1, 9)    <= sub_wire256(9);
	sub_wire2(1, 10)    <= sub_wire256(10);
	sub_wire2(1, 11)    <= sub_wire256(11);
	sub_wire2(1, 12)    <= sub_wire256(12);
	sub_wire2(1, 13)    <= sub_wire256(13);
	sub_wire2(1, 14)    <= sub_wire256(14);
	sub_wire2(1, 15)    <= sub_wire256(15);
	sub_wire2(1, 16)    <= sub_wire256(16);
	sub_wire2(1, 17)    <= sub_wire256(17);
	sub_wire2(1, 18)    <= sub_wire256(18);
	sub_wire2(1, 19)    <= sub_wire256(19);
	sub_wire2(1, 20)    <= sub_wire256(20);
	sub_wire2(1, 21)    <= sub_wire256(21);
	sub_wire2(1, 22)    <= sub_wire256(22);
	sub_wire2(1, 23)    <= sub_wire256(23);
	sub_wire2(1, 24)    <= sub_wire256(24);
	sub_wire2(1, 25)    <= sub_wire256(25);
	sub_wire2(1, 26)    <= sub_wire256(26);
	sub_wire2(1, 27)    <= sub_wire256(27);
	sub_wire2(1, 28)    <= sub_wire256(28);
	sub_wire2(1, 29)    <= sub_wire256(29);
	sub_wire2(1, 30)    <= sub_wire256(30);
	sub_wire2(1, 31)    <= sub_wire256(31);
	sub_wire2(1, 32)    <= sub_wire256(32);
	sub_wire2(1, 33)    <= sub_wire256(33);
	sub_wire2(1, 34)    <= sub_wire256(34);
	sub_wire2(1, 35)    <= sub_wire256(35);
	sub_wire2(1, 36)    <= sub_wire256(36);
	sub_wire2(1, 37)    <= sub_wire256(37);
	sub_wire2(1, 38)    <= sub_wire256(38);
	sub_wire2(1, 39)    <= sub_wire256(39);
	sub_wire2(0, 0)    <= sub_wire257(0);
	sub_wire2(0, 1)    <= sub_wire257(1);
	sub_wire2(0, 2)    <= sub_wire257(2);
	sub_wire2(0, 3)    <= sub_wire257(3);
	sub_wire2(0, 4)    <= sub_wire257(4);
	sub_wire2(0, 5)    <= sub_wire257(5);
	sub_wire2(0, 6)    <= sub_wire257(6);
	sub_wire2(0, 7)    <= sub_wire257(7);
	sub_wire2(0, 8)    <= sub_wire257(8);
	sub_wire2(0, 9)    <= sub_wire257(9);
	sub_wire2(0, 10)    <= sub_wire257(10);
	sub_wire2(0, 11)    <= sub_wire257(11);
	sub_wire2(0, 12)    <= sub_wire257(12);
	sub_wire2(0, 13)    <= sub_wire257(13);
	sub_wire2(0, 14)    <= sub_wire257(14);
	sub_wire2(0, 15)    <= sub_wire257(15);
	sub_wire2(0, 16)    <= sub_wire257(16);
	sub_wire2(0, 17)    <= sub_wire257(17);
	sub_wire2(0, 18)    <= sub_wire257(18);
	sub_wire2(0, 19)    <= sub_wire257(19);
	sub_wire2(0, 20)    <= sub_wire257(20);
	sub_wire2(0, 21)    <= sub_wire257(21);
	sub_wire2(0, 22)    <= sub_wire257(22);
	sub_wire2(0, 23)    <= sub_wire257(23);
	sub_wire2(0, 24)    <= sub_wire257(24);
	sub_wire2(0, 25)    <= sub_wire257(25);
	sub_wire2(0, 26)    <= sub_wire257(26);
	sub_wire2(0, 27)    <= sub_wire257(27);
	sub_wire2(0, 28)    <= sub_wire257(28);
	sub_wire2(0, 29)    <= sub_wire257(29);
	sub_wire2(0, 30)    <= sub_wire257(30);
	sub_wire2(0, 31)    <= sub_wire257(31);
	sub_wire2(0, 32)    <= sub_wire257(32);
	sub_wire2(0, 33)    <= sub_wire257(33);
	sub_wire2(0, 34)    <= sub_wire257(34);
	sub_wire2(0, 35)    <= sub_wire257(35);
	sub_wire2(0, 36)    <= sub_wire257(36);
	sub_wire2(0, 37)    <= sub_wire257(37);
	sub_wire2(0, 38)    <= sub_wire257(38);
	sub_wire2(0, 39)    <= sub_wire257(39);

	lpm_mux_component : lpm_mux
	GENERIC MAP (
		lpm_pipeline => 1,
		lpm_size => 256,
		lpm_type => "LPM_MUX",
		lpm_width => 40,
		lpm_widths => 8
	)
	PORT MAP (
		sel => sel,
		clock => clock,
		data => sub_wire2,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "1"
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "256"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "40"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "8"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
-- Retrieval info: USED_PORT: data0x 0 0 40 0 INPUT NODEFVAL data0x[39..0]
-- Retrieval info: USED_PORT: data100x 0 0 40 0 INPUT NODEFVAL data100x[39..0]
-- Retrieval info: USED_PORT: data101x 0 0 40 0 INPUT NODEFVAL data101x[39..0]
-- Retrieval info: USED_PORT: data102x 0 0 40 0 INPUT NODEFVAL data102x[39..0]
-- Retrieval info: USED_PORT: data103x 0 0 40 0 INPUT NODEFVAL data103x[39..0]
-- Retrieval info: USED_PORT: data104x 0 0 40 0 INPUT NODEFVAL data104x[39..0]
-- Retrieval info: USED_PORT: data105x 0 0 40 0 INPUT NODEFVAL data105x[39..0]
-- Retrieval info: USED_PORT: data106x 0 0 40 0 INPUT NODEFVAL data106x[39..0]
-- Retrieval info: USED_PORT: data107x 0 0 40 0 INPUT NODEFVAL data107x[39..0]
-- Retrieval info: USED_PORT: data108x 0 0 40 0 INPUT NODEFVAL data108x[39..0]
-- Retrieval info: USED_PORT: data109x 0 0 40 0 INPUT NODEFVAL data109x[39..0]
-- Retrieval info: USED_PORT: data10x 0 0 40 0 INPUT NODEFVAL data10x[39..0]
-- Retrieval info: USED_PORT: data110x 0 0 40 0 INPUT NODEFVAL data110x[39..0]
-- Retrieval info: USED_PORT: data111x 0 0 40 0 INPUT NODEFVAL data111x[39..0]
-- Retrieval info: USED_PORT: data112x 0 0 40 0 INPUT NODEFVAL data112x[39..0]
-- Retrieval info: USED_PORT: data113x 0 0 40 0 INPUT NODEFVAL data113x[39..0]
-- Retrieval info: USED_PORT: data114x 0 0 40 0 INPUT NODEFVAL data114x[39..0]
-- Retrieval info: USED_PORT: data115x 0 0 40 0 INPUT NODEFVAL data115x[39..0]
-- Retrieval info: USED_PORT: data116x 0 0 40 0 INPUT NODEFVAL data116x[39..0]
-- Retrieval info: USED_PORT: data117x 0 0 40 0 INPUT NODEFVAL data117x[39..0]
-- Retrieval info: USED_PORT: data118x 0 0 40 0 INPUT NODEFVAL data118x[39..0]
-- Retrieval info: USED_PORT: data119x 0 0 40 0 INPUT NODEFVAL data119x[39..0]
-- Retrieval info: USED_PORT: data11x 0 0 40 0 INPUT NODEFVAL data11x[39..0]
-- Retrieval info: USED_PORT: data120x 0 0 40 0 INPUT NODEFVAL data120x[39..0]
-- Retrieval info: USED_PORT: data121x 0 0 40 0 INPUT NODEFVAL data121x[39..0]
-- Retrieval info: USED_PORT: data122x 0 0 40 0 INPUT NODEFVAL data122x[39..0]
-- Retrieval info: USED_PORT: data123x 0 0 40 0 INPUT NODEFVAL data123x[39..0]
-- Retrieval info: USED_PORT: data124x 0 0 40 0 INPUT NODEFVAL data124x[39..0]
-- Retrieval info: USED_PORT: data125x 0 0 40 0 INPUT NODEFVAL data125x[39..0]
-- Retrieval info: USED_PORT: data126x 0 0 40 0 INPUT NODEFVAL data126x[39..0]
-- Retrieval info: USED_PORT: data127x 0 0 40 0 INPUT NODEFVAL data127x[39..0]
-- Retrieval info: USED_PORT: data128x 0 0 40 0 INPUT NODEFVAL data128x[39..0]
-- Retrieval info: USED_PORT: data129x 0 0 40 0 INPUT NODEFVAL data129x[39..0]
-- Retrieval info: USED_PORT: data12x 0 0 40 0 INPUT NODEFVAL data12x[39..0]
-- Retrieval info: USED_PORT: data130x 0 0 40 0 INPUT NODEFVAL data130x[39..0]
-- Retrieval info: USED_PORT: data131x 0 0 40 0 INPUT NODEFVAL data131x[39..0]
-- Retrieval info: USED_PORT: data132x 0 0 40 0 INPUT NODEFVAL data132x[39..0]
-- Retrieval info: USED_PORT: data133x 0 0 40 0 INPUT NODEFVAL data133x[39..0]
-- Retrieval info: USED_PORT: data134x 0 0 40 0 INPUT NODEFVAL data134x[39..0]
-- Retrieval info: USED_PORT: data135x 0 0 40 0 INPUT NODEFVAL data135x[39..0]
-- Retrieval info: USED_PORT: data136x 0 0 40 0 INPUT NODEFVAL data136x[39..0]
-- Retrieval info: USED_PORT: data137x 0 0 40 0 INPUT NODEFVAL data137x[39..0]
-- Retrieval info: USED_PORT: data138x 0 0 40 0 INPUT NODEFVAL data138x[39..0]
-- Retrieval info: USED_PORT: data139x 0 0 40 0 INPUT NODEFVAL data139x[39..0]
-- Retrieval info: USED_PORT: data13x 0 0 40 0 INPUT NODEFVAL data13x[39..0]
-- Retrieval info: USED_PORT: data140x 0 0 40 0 INPUT NODEFVAL data140x[39..0]
-- Retrieval info: USED_PORT: data141x 0 0 40 0 INPUT NODEFVAL data141x[39..0]
-- Retrieval info: USED_PORT: data142x 0 0 40 0 INPUT NODEFVAL data142x[39..0]
-- Retrieval info: USED_PORT: data143x 0 0 40 0 INPUT NODEFVAL data143x[39..0]
-- Retrieval info: USED_PORT: data144x 0 0 40 0 INPUT NODEFVAL data144x[39..0]
-- Retrieval info: USED_PORT: data145x 0 0 40 0 INPUT NODEFVAL data145x[39..0]
-- Retrieval info: USED_PORT: data146x 0 0 40 0 INPUT NODEFVAL data146x[39..0]
-- Retrieval info: USED_PORT: data147x 0 0 40 0 INPUT NODEFVAL data147x[39..0]
-- Retrieval info: USED_PORT: data148x 0 0 40 0 INPUT NODEFVAL data148x[39..0]
-- Retrieval info: USED_PORT: data149x 0 0 40 0 INPUT NODEFVAL data149x[39..0]
-- Retrieval info: USED_PORT: data14x 0 0 40 0 INPUT NODEFVAL data14x[39..0]
-- Retrieval info: USED_PORT: data150x 0 0 40 0 INPUT NODEFVAL data150x[39..0]
-- Retrieval info: USED_PORT: data151x 0 0 40 0 INPUT NODEFVAL data151x[39..0]
-- Retrieval info: USED_PORT: data152x 0 0 40 0 INPUT NODEFVAL data152x[39..0]
-- Retrieval info: USED_PORT: data153x 0 0 40 0 INPUT NODEFVAL data153x[39..0]
-- Retrieval info: USED_PORT: data154x 0 0 40 0 INPUT NODEFVAL data154x[39..0]
-- Retrieval info: USED_PORT: data155x 0 0 40 0 INPUT NODEFVAL data155x[39..0]
-- Retrieval info: USED_PORT: data156x 0 0 40 0 INPUT NODEFVAL data156x[39..0]
-- Retrieval info: USED_PORT: data157x 0 0 40 0 INPUT NODEFVAL data157x[39..0]
-- Retrieval info: USED_PORT: data158x 0 0 40 0 INPUT NODEFVAL data158x[39..0]
-- Retrieval info: USED_PORT: data159x 0 0 40 0 INPUT NODEFVAL data159x[39..0]
-- Retrieval info: USED_PORT: data15x 0 0 40 0 INPUT NODEFVAL data15x[39..0]
-- Retrieval info: USED_PORT: data160x 0 0 40 0 INPUT NODEFVAL data160x[39..0]
-- Retrieval info: USED_PORT: data161x 0 0 40 0 INPUT NODEFVAL data161x[39..0]
-- Retrieval info: USED_PORT: data162x 0 0 40 0 INPUT NODEFVAL data162x[39..0]
-- Retrieval info: USED_PORT: data163x 0 0 40 0 INPUT NODEFVAL data163x[39..0]
-- Retrieval info: USED_PORT: data164x 0 0 40 0 INPUT NODEFVAL data164x[39..0]
-- Retrieval info: USED_PORT: data165x 0 0 40 0 INPUT NODEFVAL data165x[39..0]
-- Retrieval info: USED_PORT: data166x 0 0 40 0 INPUT NODEFVAL data166x[39..0]
-- Retrieval info: USED_PORT: data167x 0 0 40 0 INPUT NODEFVAL data167x[39..0]
-- Retrieval info: USED_PORT: data168x 0 0 40 0 INPUT NODEFVAL data168x[39..0]
-- Retrieval info: USED_PORT: data169x 0 0 40 0 INPUT NODEFVAL data169x[39..0]
-- Retrieval info: USED_PORT: data16x 0 0 40 0 INPUT NODEFVAL data16x[39..0]
-- Retrieval info: USED_PORT: data170x 0 0 40 0 INPUT NODEFVAL data170x[39..0]
-- Retrieval info: USED_PORT: data171x 0 0 40 0 INPUT NODEFVAL data171x[39..0]
-- Retrieval info: USED_PORT: data172x 0 0 40 0 INPUT NODEFVAL data172x[39..0]
-- Retrieval info: USED_PORT: data173x 0 0 40 0 INPUT NODEFVAL data173x[39..0]
-- Retrieval info: USED_PORT: data174x 0 0 40 0 INPUT NODEFVAL data174x[39..0]
-- Retrieval info: USED_PORT: data175x 0 0 40 0 INPUT NODEFVAL data175x[39..0]
-- Retrieval info: USED_PORT: data176x 0 0 40 0 INPUT NODEFVAL data176x[39..0]
-- Retrieval info: USED_PORT: data177x 0 0 40 0 INPUT NODEFVAL data177x[39..0]
-- Retrieval info: USED_PORT: data178x 0 0 40 0 INPUT NODEFVAL data178x[39..0]
-- Retrieval info: USED_PORT: data179x 0 0 40 0 INPUT NODEFVAL data179x[39..0]
-- Retrieval info: USED_PORT: data17x 0 0 40 0 INPUT NODEFVAL data17x[39..0]
-- Retrieval info: USED_PORT: data180x 0 0 40 0 INPUT NODEFVAL data180x[39..0]
-- Retrieval info: USED_PORT: data181x 0 0 40 0 INPUT NODEFVAL data181x[39..0]
-- Retrieval info: USED_PORT: data182x 0 0 40 0 INPUT NODEFVAL data182x[39..0]
-- Retrieval info: USED_PORT: data183x 0 0 40 0 INPUT NODEFVAL data183x[39..0]
-- Retrieval info: USED_PORT: data184x 0 0 40 0 INPUT NODEFVAL data184x[39..0]
-- Retrieval info: USED_PORT: data185x 0 0 40 0 INPUT NODEFVAL data185x[39..0]
-- Retrieval info: USED_PORT: data186x 0 0 40 0 INPUT NODEFVAL data186x[39..0]
-- Retrieval info: USED_PORT: data187x 0 0 40 0 INPUT NODEFVAL data187x[39..0]
-- Retrieval info: USED_PORT: data188x 0 0 40 0 INPUT NODEFVAL data188x[39..0]
-- Retrieval info: USED_PORT: data189x 0 0 40 0 INPUT NODEFVAL data189x[39..0]
-- Retrieval info: USED_PORT: data18x 0 0 40 0 INPUT NODEFVAL data18x[39..0]
-- Retrieval info: USED_PORT: data190x 0 0 40 0 INPUT NODEFVAL data190x[39..0]
-- Retrieval info: USED_PORT: data191x 0 0 40 0 INPUT NODEFVAL data191x[39..0]
-- Retrieval info: USED_PORT: data192x 0 0 40 0 INPUT NODEFVAL data192x[39..0]
-- Retrieval info: USED_PORT: data193x 0 0 40 0 INPUT NODEFVAL data193x[39..0]
-- Retrieval info: USED_PORT: data194x 0 0 40 0 INPUT NODEFVAL data194x[39..0]
-- Retrieval info: USED_PORT: data195x 0 0 40 0 INPUT NODEFVAL data195x[39..0]
-- Retrieval info: USED_PORT: data196x 0 0 40 0 INPUT NODEFVAL data196x[39..0]
-- Retrieval info: USED_PORT: data197x 0 0 40 0 INPUT NODEFVAL data197x[39..0]
-- Retrieval info: USED_PORT: data198x 0 0 40 0 INPUT NODEFVAL data198x[39..0]
-- Retrieval info: USED_PORT: data199x 0 0 40 0 INPUT NODEFVAL data199x[39..0]
-- Retrieval info: USED_PORT: data19x 0 0 40 0 INPUT NODEFVAL data19x[39..0]
-- Retrieval info: USED_PORT: data1x 0 0 40 0 INPUT NODEFVAL data1x[39..0]
-- Retrieval info: USED_PORT: data200x 0 0 40 0 INPUT NODEFVAL data200x[39..0]
-- Retrieval info: USED_PORT: data201x 0 0 40 0 INPUT NODEFVAL data201x[39..0]
-- Retrieval info: USED_PORT: data202x 0 0 40 0 INPUT NODEFVAL data202x[39..0]
-- Retrieval info: USED_PORT: data203x 0 0 40 0 INPUT NODEFVAL data203x[39..0]
-- Retrieval info: USED_PORT: data204x 0 0 40 0 INPUT NODEFVAL data204x[39..0]
-- Retrieval info: USED_PORT: data205x 0 0 40 0 INPUT NODEFVAL data205x[39..0]
-- Retrieval info: USED_PORT: data206x 0 0 40 0 INPUT NODEFVAL data206x[39..0]
-- Retrieval info: USED_PORT: data207x 0 0 40 0 INPUT NODEFVAL data207x[39..0]
-- Retrieval info: USED_PORT: data208x 0 0 40 0 INPUT NODEFVAL data208x[39..0]
-- Retrieval info: USED_PORT: data209x 0 0 40 0 INPUT NODEFVAL data209x[39..0]
-- Retrieval info: USED_PORT: data20x 0 0 40 0 INPUT NODEFVAL data20x[39..0]
-- Retrieval info: USED_PORT: data210x 0 0 40 0 INPUT NODEFVAL data210x[39..0]
-- Retrieval info: USED_PORT: data211x 0 0 40 0 INPUT NODEFVAL data211x[39..0]
-- Retrieval info: USED_PORT: data212x 0 0 40 0 INPUT NODEFVAL data212x[39..0]
-- Retrieval info: USED_PORT: data213x 0 0 40 0 INPUT NODEFVAL data213x[39..0]
-- Retrieval info: USED_PORT: data214x 0 0 40 0 INPUT NODEFVAL data214x[39..0]
-- Retrieval info: USED_PORT: data215x 0 0 40 0 INPUT NODEFVAL data215x[39..0]
-- Retrieval info: USED_PORT: data216x 0 0 40 0 INPUT NODEFVAL data216x[39..0]
-- Retrieval info: USED_PORT: data217x 0 0 40 0 INPUT NODEFVAL data217x[39..0]
-- Retrieval info: USED_PORT: data218x 0 0 40 0 INPUT NODEFVAL data218x[39..0]
-- Retrieval info: USED_PORT: data219x 0 0 40 0 INPUT NODEFVAL data219x[39..0]
-- Retrieval info: USED_PORT: data21x 0 0 40 0 INPUT NODEFVAL data21x[39..0]
-- Retrieval info: USED_PORT: data220x 0 0 40 0 INPUT NODEFVAL data220x[39..0]
-- Retrieval info: USED_PORT: data221x 0 0 40 0 INPUT NODEFVAL data221x[39..0]
-- Retrieval info: USED_PORT: data222x 0 0 40 0 INPUT NODEFVAL data222x[39..0]
-- Retrieval info: USED_PORT: data223x 0 0 40 0 INPUT NODEFVAL data223x[39..0]
-- Retrieval info: USED_PORT: data224x 0 0 40 0 INPUT NODEFVAL data224x[39..0]
-- Retrieval info: USED_PORT: data225x 0 0 40 0 INPUT NODEFVAL data225x[39..0]
-- Retrieval info: USED_PORT: data226x 0 0 40 0 INPUT NODEFVAL data226x[39..0]
-- Retrieval info: USED_PORT: data227x 0 0 40 0 INPUT NODEFVAL data227x[39..0]
-- Retrieval info: USED_PORT: data228x 0 0 40 0 INPUT NODEFVAL data228x[39..0]
-- Retrieval info: USED_PORT: data229x 0 0 40 0 INPUT NODEFVAL data229x[39..0]
-- Retrieval info: USED_PORT: data22x 0 0 40 0 INPUT NODEFVAL data22x[39..0]
-- Retrieval info: USED_PORT: data230x 0 0 40 0 INPUT NODEFVAL data230x[39..0]
-- Retrieval info: USED_PORT: data231x 0 0 40 0 INPUT NODEFVAL data231x[39..0]
-- Retrieval info: USED_PORT: data232x 0 0 40 0 INPUT NODEFVAL data232x[39..0]
-- Retrieval info: USED_PORT: data233x 0 0 40 0 INPUT NODEFVAL data233x[39..0]
-- Retrieval info: USED_PORT: data234x 0 0 40 0 INPUT NODEFVAL data234x[39..0]
-- Retrieval info: USED_PORT: data235x 0 0 40 0 INPUT NODEFVAL data235x[39..0]
-- Retrieval info: USED_PORT: data236x 0 0 40 0 INPUT NODEFVAL data236x[39..0]
-- Retrieval info: USED_PORT: data237x 0 0 40 0 INPUT NODEFVAL data237x[39..0]
-- Retrieval info: USED_PORT: data238x 0 0 40 0 INPUT NODEFVAL data238x[39..0]
-- Retrieval info: USED_PORT: data239x 0 0 40 0 INPUT NODEFVAL data239x[39..0]
-- Retrieval info: USED_PORT: data23x 0 0 40 0 INPUT NODEFVAL data23x[39..0]
-- Retrieval info: USED_PORT: data240x 0 0 40 0 INPUT NODEFVAL data240x[39..0]
-- Retrieval info: USED_PORT: data241x 0 0 40 0 INPUT NODEFVAL data241x[39..0]
-- Retrieval info: USED_PORT: data242x 0 0 40 0 INPUT NODEFVAL data242x[39..0]
-- Retrieval info: USED_PORT: data243x 0 0 40 0 INPUT NODEFVAL data243x[39..0]
-- Retrieval info: USED_PORT: data244x 0 0 40 0 INPUT NODEFVAL data244x[39..0]
-- Retrieval info: USED_PORT: data245x 0 0 40 0 INPUT NODEFVAL data245x[39..0]
-- Retrieval info: USED_PORT: data246x 0 0 40 0 INPUT NODEFVAL data246x[39..0]
-- Retrieval info: USED_PORT: data247x 0 0 40 0 INPUT NODEFVAL data247x[39..0]
-- Retrieval info: USED_PORT: data248x 0 0 40 0 INPUT NODEFVAL data248x[39..0]
-- Retrieval info: USED_PORT: data249x 0 0 40 0 INPUT NODEFVAL data249x[39..0]
-- Retrieval info: USED_PORT: data24x 0 0 40 0 INPUT NODEFVAL data24x[39..0]
-- Retrieval info: USED_PORT: data250x 0 0 40 0 INPUT NODEFVAL data250x[39..0]
-- Retrieval info: USED_PORT: data251x 0 0 40 0 INPUT NODEFVAL data251x[39..0]
-- Retrieval info: USED_PORT: data252x 0 0 40 0 INPUT NODEFVAL data252x[39..0]
-- Retrieval info: USED_PORT: data253x 0 0 40 0 INPUT NODEFVAL data253x[39..0]
-- Retrieval info: USED_PORT: data254x 0 0 40 0 INPUT NODEFVAL data254x[39..0]
-- Retrieval info: USED_PORT: data255x 0 0 40 0 INPUT NODEFVAL data255x[39..0]
-- Retrieval info: USED_PORT: data25x 0 0 40 0 INPUT NODEFVAL data25x[39..0]
-- Retrieval info: USED_PORT: data26x 0 0 40 0 INPUT NODEFVAL data26x[39..0]
-- Retrieval info: USED_PORT: data27x 0 0 40 0 INPUT NODEFVAL data27x[39..0]
-- Retrieval info: USED_PORT: data28x 0 0 40 0 INPUT NODEFVAL data28x[39..0]
-- Retrieval info: USED_PORT: data29x 0 0 40 0 INPUT NODEFVAL data29x[39..0]
-- Retrieval info: USED_PORT: data2x 0 0 40 0 INPUT NODEFVAL data2x[39..0]
-- Retrieval info: USED_PORT: data30x 0 0 40 0 INPUT NODEFVAL data30x[39..0]
-- Retrieval info: USED_PORT: data31x 0 0 40 0 INPUT NODEFVAL data31x[39..0]
-- Retrieval info: USED_PORT: data32x 0 0 40 0 INPUT NODEFVAL data32x[39..0]
-- Retrieval info: USED_PORT: data33x 0 0 40 0 INPUT NODEFVAL data33x[39..0]
-- Retrieval info: USED_PORT: data34x 0 0 40 0 INPUT NODEFVAL data34x[39..0]
-- Retrieval info: USED_PORT: data35x 0 0 40 0 INPUT NODEFVAL data35x[39..0]
-- Retrieval info: USED_PORT: data36x 0 0 40 0 INPUT NODEFVAL data36x[39..0]
-- Retrieval info: USED_PORT: data37x 0 0 40 0 INPUT NODEFVAL data37x[39..0]
-- Retrieval info: USED_PORT: data38x 0 0 40 0 INPUT NODEFVAL data38x[39..0]
-- Retrieval info: USED_PORT: data39x 0 0 40 0 INPUT NODEFVAL data39x[39..0]
-- Retrieval info: USED_PORT: data3x 0 0 40 0 INPUT NODEFVAL data3x[39..0]
-- Retrieval info: USED_PORT: data40x 0 0 40 0 INPUT NODEFVAL data40x[39..0]
-- Retrieval info: USED_PORT: data41x 0 0 40 0 INPUT NODEFVAL data41x[39..0]
-- Retrieval info: USED_PORT: data42x 0 0 40 0 INPUT NODEFVAL data42x[39..0]
-- Retrieval info: USED_PORT: data43x 0 0 40 0 INPUT NODEFVAL data43x[39..0]
-- Retrieval info: USED_PORT: data44x 0 0 40 0 INPUT NODEFVAL data44x[39..0]
-- Retrieval info: USED_PORT: data45x 0 0 40 0 INPUT NODEFVAL data45x[39..0]
-- Retrieval info: USED_PORT: data46x 0 0 40 0 INPUT NODEFVAL data46x[39..0]
-- Retrieval info: USED_PORT: data47x 0 0 40 0 INPUT NODEFVAL data47x[39..0]
-- Retrieval info: USED_PORT: data48x 0 0 40 0 INPUT NODEFVAL data48x[39..0]
-- Retrieval info: USED_PORT: data49x 0 0 40 0 INPUT NODEFVAL data49x[39..0]
-- Retrieval info: USED_PORT: data4x 0 0 40 0 INPUT NODEFVAL data4x[39..0]
-- Retrieval info: USED_PORT: data50x 0 0 40 0 INPUT NODEFVAL data50x[39..0]
-- Retrieval info: USED_PORT: data51x 0 0 40 0 INPUT NODEFVAL data51x[39..0]
-- Retrieval info: USED_PORT: data52x 0 0 40 0 INPUT NODEFVAL data52x[39..0]
-- Retrieval info: USED_PORT: data53x 0 0 40 0 INPUT NODEFVAL data53x[39..0]
-- Retrieval info: USED_PORT: data54x 0 0 40 0 INPUT NODEFVAL data54x[39..0]
-- Retrieval info: USED_PORT: data55x 0 0 40 0 INPUT NODEFVAL data55x[39..0]
-- Retrieval info: USED_PORT: data56x 0 0 40 0 INPUT NODEFVAL data56x[39..0]
-- Retrieval info: USED_PORT: data57x 0 0 40 0 INPUT NODEFVAL data57x[39..0]
-- Retrieval info: USED_PORT: data58x 0 0 40 0 INPUT NODEFVAL data58x[39..0]
-- Retrieval info: USED_PORT: data59x 0 0 40 0 INPUT NODEFVAL data59x[39..0]
-- Retrieval info: USED_PORT: data5x 0 0 40 0 INPUT NODEFVAL data5x[39..0]
-- Retrieval info: USED_PORT: data60x 0 0 40 0 INPUT NODEFVAL data60x[39..0]
-- Retrieval info: USED_PORT: data61x 0 0 40 0 INPUT NODEFVAL data61x[39..0]
-- Retrieval info: USED_PORT: data62x 0 0 40 0 INPUT NODEFVAL data62x[39..0]
-- Retrieval info: USED_PORT: data63x 0 0 40 0 INPUT NODEFVAL data63x[39..0]
-- Retrieval info: USED_PORT: data64x 0 0 40 0 INPUT NODEFVAL data64x[39..0]
-- Retrieval info: USED_PORT: data65x 0 0 40 0 INPUT NODEFVAL data65x[39..0]
-- Retrieval info: USED_PORT: data66x 0 0 40 0 INPUT NODEFVAL data66x[39..0]
-- Retrieval info: USED_PORT: data67x 0 0 40 0 INPUT NODEFVAL data67x[39..0]
-- Retrieval info: USED_PORT: data68x 0 0 40 0 INPUT NODEFVAL data68x[39..0]
-- Retrieval info: USED_PORT: data69x 0 0 40 0 INPUT NODEFVAL data69x[39..0]
-- Retrieval info: USED_PORT: data6x 0 0 40 0 INPUT NODEFVAL data6x[39..0]
-- Retrieval info: USED_PORT: data70x 0 0 40 0 INPUT NODEFVAL data70x[39..0]
-- Retrieval info: USED_PORT: data71x 0 0 40 0 INPUT NODEFVAL data71x[39..0]
-- Retrieval info: USED_PORT: data72x 0 0 40 0 INPUT NODEFVAL data72x[39..0]
-- Retrieval info: USED_PORT: data73x 0 0 40 0 INPUT NODEFVAL data73x[39..0]
-- Retrieval info: USED_PORT: data74x 0 0 40 0 INPUT NODEFVAL data74x[39..0]
-- Retrieval info: USED_PORT: data75x 0 0 40 0 INPUT NODEFVAL data75x[39..0]
-- Retrieval info: USED_PORT: data76x 0 0 40 0 INPUT NODEFVAL data76x[39..0]
-- Retrieval info: USED_PORT: data77x 0 0 40 0 INPUT NODEFVAL data77x[39..0]
-- Retrieval info: USED_PORT: data78x 0 0 40 0 INPUT NODEFVAL data78x[39..0]
-- Retrieval info: USED_PORT: data79x 0 0 40 0 INPUT NODEFVAL data79x[39..0]
-- Retrieval info: USED_PORT: data7x 0 0 40 0 INPUT NODEFVAL data7x[39..0]
-- Retrieval info: USED_PORT: data80x 0 0 40 0 INPUT NODEFVAL data80x[39..0]
-- Retrieval info: USED_PORT: data81x 0 0 40 0 INPUT NODEFVAL data81x[39..0]
-- Retrieval info: USED_PORT: data82x 0 0 40 0 INPUT NODEFVAL data82x[39..0]
-- Retrieval info: USED_PORT: data83x 0 0 40 0 INPUT NODEFVAL data83x[39..0]
-- Retrieval info: USED_PORT: data84x 0 0 40 0 INPUT NODEFVAL data84x[39..0]
-- Retrieval info: USED_PORT: data85x 0 0 40 0 INPUT NODEFVAL data85x[39..0]
-- Retrieval info: USED_PORT: data86x 0 0 40 0 INPUT NODEFVAL data86x[39..0]
-- Retrieval info: USED_PORT: data87x 0 0 40 0 INPUT NODEFVAL data87x[39..0]
-- Retrieval info: USED_PORT: data88x 0 0 40 0 INPUT NODEFVAL data88x[39..0]
-- Retrieval info: USED_PORT: data89x 0 0 40 0 INPUT NODEFVAL data89x[39..0]
-- Retrieval info: USED_PORT: data8x 0 0 40 0 INPUT NODEFVAL data8x[39..0]
-- Retrieval info: USED_PORT: data90x 0 0 40 0 INPUT NODEFVAL data90x[39..0]
-- Retrieval info: USED_PORT: data91x 0 0 40 0 INPUT NODEFVAL data91x[39..0]
-- Retrieval info: USED_PORT: data92x 0 0 40 0 INPUT NODEFVAL data92x[39..0]
-- Retrieval info: USED_PORT: data93x 0 0 40 0 INPUT NODEFVAL data93x[39..0]
-- Retrieval info: USED_PORT: data94x 0 0 40 0 INPUT NODEFVAL data94x[39..0]
-- Retrieval info: USED_PORT: data95x 0 0 40 0 INPUT NODEFVAL data95x[39..0]
-- Retrieval info: USED_PORT: data96x 0 0 40 0 INPUT NODEFVAL data96x[39..0]
-- Retrieval info: USED_PORT: data97x 0 0 40 0 INPUT NODEFVAL data97x[39..0]
-- Retrieval info: USED_PORT: data98x 0 0 40 0 INPUT NODEFVAL data98x[39..0]
-- Retrieval info: USED_PORT: data99x 0 0 40 0 INPUT NODEFVAL data99x[39..0]
-- Retrieval info: USED_PORT: data9x 0 0 40 0 INPUT NODEFVAL data9x[39..0]
-- Retrieval info: USED_PORT: result 0 0 40 0 OUTPUT NODEFVAL result[39..0]
-- Retrieval info: USED_PORT: sel 0 0 8 0 INPUT NODEFVAL sel[7..0]
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: result 0 0 40 0 @result 0 0 40 0
-- Retrieval info: CONNECT: @data 1 255 40 0 data255x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 254 40 0 data254x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 253 40 0 data253x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 252 40 0 data252x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 251 40 0 data251x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 250 40 0 data250x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 249 40 0 data249x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 248 40 0 data248x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 247 40 0 data247x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 246 40 0 data246x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 245 40 0 data245x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 244 40 0 data244x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 243 40 0 data243x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 242 40 0 data242x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 241 40 0 data241x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 240 40 0 data240x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 239 40 0 data239x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 238 40 0 data238x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 237 40 0 data237x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 236 40 0 data236x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 235 40 0 data235x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 234 40 0 data234x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 233 40 0 data233x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 232 40 0 data232x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 231 40 0 data231x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 230 40 0 data230x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 229 40 0 data229x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 228 40 0 data228x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 227 40 0 data227x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 226 40 0 data226x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 225 40 0 data225x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 224 40 0 data224x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 223 40 0 data223x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 222 40 0 data222x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 221 40 0 data221x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 220 40 0 data220x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 219 40 0 data219x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 218 40 0 data218x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 217 40 0 data217x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 216 40 0 data216x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 215 40 0 data215x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 214 40 0 data214x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 213 40 0 data213x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 212 40 0 data212x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 211 40 0 data211x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 210 40 0 data210x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 209 40 0 data209x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 208 40 0 data208x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 207 40 0 data207x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 206 40 0 data206x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 205 40 0 data205x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 204 40 0 data204x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 203 40 0 data203x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 202 40 0 data202x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 201 40 0 data201x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 200 40 0 data200x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 199 40 0 data199x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 198 40 0 data198x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 197 40 0 data197x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 196 40 0 data196x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 195 40 0 data195x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 194 40 0 data194x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 193 40 0 data193x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 192 40 0 data192x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 191 40 0 data191x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 190 40 0 data190x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 189 40 0 data189x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 188 40 0 data188x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 187 40 0 data187x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 186 40 0 data186x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 185 40 0 data185x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 184 40 0 data184x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 183 40 0 data183x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 182 40 0 data182x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 181 40 0 data181x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 180 40 0 data180x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 179 40 0 data179x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 178 40 0 data178x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 177 40 0 data177x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 176 40 0 data176x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 175 40 0 data175x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 174 40 0 data174x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 173 40 0 data173x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 172 40 0 data172x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 171 40 0 data171x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 170 40 0 data170x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 169 40 0 data169x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 168 40 0 data168x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 167 40 0 data167x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 166 40 0 data166x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 165 40 0 data165x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 164 40 0 data164x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 163 40 0 data163x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 162 40 0 data162x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 161 40 0 data161x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 160 40 0 data160x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 159 40 0 data159x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 158 40 0 data158x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 157 40 0 data157x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 156 40 0 data156x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 155 40 0 data155x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 154 40 0 data154x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 153 40 0 data153x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 152 40 0 data152x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 151 40 0 data151x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 150 40 0 data150x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 149 40 0 data149x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 148 40 0 data148x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 147 40 0 data147x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 146 40 0 data146x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 145 40 0 data145x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 144 40 0 data144x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 143 40 0 data143x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 142 40 0 data142x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 141 40 0 data141x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 140 40 0 data140x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 139 40 0 data139x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 138 40 0 data138x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 137 40 0 data137x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 136 40 0 data136x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 135 40 0 data135x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 134 40 0 data134x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 133 40 0 data133x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 132 40 0 data132x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 131 40 0 data131x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 130 40 0 data130x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 129 40 0 data129x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 128 40 0 data128x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 127 40 0 data127x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 126 40 0 data126x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 125 40 0 data125x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 124 40 0 data124x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 123 40 0 data123x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 122 40 0 data122x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 121 40 0 data121x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 120 40 0 data120x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 119 40 0 data119x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 118 40 0 data118x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 117 40 0 data117x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 116 40 0 data116x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 115 40 0 data115x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 114 40 0 data114x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 113 40 0 data113x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 112 40 0 data112x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 111 40 0 data111x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 110 40 0 data110x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 109 40 0 data109x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 108 40 0 data108x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 107 40 0 data107x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 106 40 0 data106x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 105 40 0 data105x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 104 40 0 data104x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 103 40 0 data103x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 102 40 0 data102x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 101 40 0 data101x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 100 40 0 data100x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 99 40 0 data99x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 98 40 0 data98x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 97 40 0 data97x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 96 40 0 data96x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 95 40 0 data95x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 94 40 0 data94x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 93 40 0 data93x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 92 40 0 data92x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 91 40 0 data91x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 90 40 0 data90x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 89 40 0 data89x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 88 40 0 data88x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 87 40 0 data87x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 86 40 0 data86x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 85 40 0 data85x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 84 40 0 data84x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 83 40 0 data83x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 82 40 0 data82x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 81 40 0 data81x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 80 40 0 data80x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 79 40 0 data79x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 78 40 0 data78x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 77 40 0 data77x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 76 40 0 data76x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 75 40 0 data75x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 74 40 0 data74x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 73 40 0 data73x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 72 40 0 data72x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 71 40 0 data71x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 70 40 0 data70x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 69 40 0 data69x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 68 40 0 data68x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 67 40 0 data67x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 66 40 0 data66x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 65 40 0 data65x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 64 40 0 data64x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 63 40 0 data63x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 62 40 0 data62x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 61 40 0 data61x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 60 40 0 data60x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 59 40 0 data59x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 58 40 0 data58x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 57 40 0 data57x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 56 40 0 data56x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 55 40 0 data55x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 54 40 0 data54x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 53 40 0 data53x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 52 40 0 data52x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 51 40 0 data51x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 50 40 0 data50x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 49 40 0 data49x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 48 40 0 data48x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 47 40 0 data47x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 46 40 0 data46x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 45 40 0 data45x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 44 40 0 data44x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 43 40 0 data43x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 42 40 0 data42x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 41 40 0 data41x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 40 40 0 data40x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 39 40 0 data39x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 38 40 0 data38x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 37 40 0 data37x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 36 40 0 data36x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 35 40 0 data35x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 34 40 0 data34x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 33 40 0 data33x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 32 40 0 data32x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 31 40 0 data31x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 30 40 0 data30x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 29 40 0 data29x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 28 40 0 data28x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 27 40 0 data27x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 26 40 0 data26x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 25 40 0 data25x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 24 40 0 data24x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 23 40 0 data23x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 22 40 0 data22x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 21 40 0 data21x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 20 40 0 data20x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 19 40 0 data19x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 18 40 0 data18x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 17 40 0 data17x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 16 40 0 data16x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 15 40 0 data15x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 14 40 0 data14x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 13 40 0 data13x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 12 40 0 data12x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 11 40 0 data11x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 10 40 0 data10x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 9 40 0 data9x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 8 40 0 data8x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 7 40 0 data7x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 6 40 0 data6x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 5 40 0 data5x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 4 40 0 data4x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 3 40 0 data3x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 2 40 0 data2x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 1 40 0 data1x 0 0 40 0
-- Retrieval info: CONNECT: @data 1 0 40 0 data0x 0 0 40 0
-- Retrieval info: CONNECT: @sel 0 0 8 0 sel 0 0 8 0
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
