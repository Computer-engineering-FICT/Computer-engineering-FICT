* /root/laba1/2.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 

*----------------------------------------------

V_V1 2 0 dc 0.0 ac 1.0 sin(0.0 10 10000 0 0) 
C_C1 1 0 0.59n IC=0 
R_R1 2 1 100000 

*----------------------------------------------

.tran 2e-06 0.0003 0 UIC
.print tran  v(2)
.op

.end
