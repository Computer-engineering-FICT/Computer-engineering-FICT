* /root/laba11/1.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/UA741.model


*----------------------------------------------

M_M1 5 12 7 0 nmos 
M_M2 7 4 6 0 nmos 
V_V1 11 0 dc 0.0 ac 0.0 sin(5 1 50000 0 0) 
V_V2 3 0 dc 0.0 ac 0.0 sin(5 1 10000 0 0) 
R_R1 3 5 5k 
R_R2 11 6 1k 
V_V3 12 0 dc 0.0 ac 0.0 PULSE 0.0 17 0.0 0.001u 0.001u 100u 200u 
V_V4 10 4 dc 0.0 ac 0.0 PULSE 0.0 17 0 0.001u 0.001u 100u 200u 
V_V5 10 0 dc 15 
V_V7 8 0 dc 5 
Q_Q1 8 1 2 NPN 
R_R4 2 9 500 
V_V6 0 9 dc 5 
R_R3 2 0 50 
.model nmos nmos (vto=3.63886 KP=20u  gamma=0 phi=600m lambda=35.07m rd=1.10826 rs=187.488m cbd=397.524p cgso=617.586p cgdo=617.586p tox=0 nsub=0 tpg=1 uo=600 ) 
X_U1 7 2 8 9 1 UA741 
.model NPN NPN (is=3.0E-14 NF=1.0 BF=200 IKF=0.5 VAF=100 ISE=7.5E-15 NE=1.4 NR=1.0 BR=4 IKR=0.24 VAR=28 ISC=1.0E-11 NC=1.4 RB=0.1 RE=0.2 RC=0.1 CJC=9.0E-12 MJC=0.35 VJC=0.4 CJE=27.0E-12 TF=0.3E-9 TR=100E-9) 

*----------------------------------------------

.tran 5e-05 0.0005 0 UIC
.print tran  v(7)
.op

.end
