*This subcircuit models the PAL16C1 from National
*
.subckt PAL16C1 1 2 3 4 5 6 7 8 9 11 12 13 14 15 16 17 18 19
+     optional:  20=$G_DPWR 10=$G_DGND
+     params:  MNTYMXDLY=0 IO_LEVEL=0
+     text: JEDFILE="PAL16C1.JED"

U1 PLANDC(16,16) 20 10
+  2 1 3 19 4 18 5 17 6 14 7 13 8 12 9 11
+  ROW1 ROW2 ROW3 ROW4 ROW5 ROW6 ROW7 ROW8 ROW9 ROW10
+  ROW11 ROW12 ROW13 ROW14 ROW15 ROW16
+  DLY_16C1 IO_LS MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}
+  FILE=|JEDFILE|

U2 ORA(8,2) 20 10
+  ROW1 ROW2 ROW3 ROW4 ROW5 ROW6 ROW7 ROW8
+  ROW9 ROW10 ROW11 ROW12 ROW13 ROW14 ROW15 ROW16
+  OR1 OR2
+  D0_GATE IO_LS MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U3 OR(2) 20 10
+  OR1 OR2 16
+  D0_GATE IO_LS MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U4 NOR(2) 20 10
+  OR1 OR2 15
+  D0_GATE IO_LS MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

.model DLY_16C1 upld (tplhTY=25ns tplhMX=35ns tphlTY=25ns tphlMX=35ns)

.ENDS

