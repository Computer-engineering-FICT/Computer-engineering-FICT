* /root/laba4/4_1.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 

*----------------------------------------------

V_V2 1 0 dc 10 
V_V1 3 0 dc 0.0 ac 0.0 sin(0.0 1 10meg 0 0) 
.model nmos nmos (vto=3.63886 KP=20u  gamma=0 phi=600m lambda=35.07m rd=1.10826 rs=187.488m cbd=397.524p cgso=617.586p cgdo=617.586p tox=0 nsub=0 tpg=1 uo=600 ) 
M_M1 2 3 0 0 nmos 
R_R1 2 1 45000 
Vtpi@1 1 2 0
*----------------------------------------------

.dc V_V1 0 5 0.1
.print dc   v(1)
.op

.end
