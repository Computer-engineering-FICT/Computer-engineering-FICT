* /root/laba7/21.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/UA741.model

*----------------------------------------------

V_V1 5 0 dc 0.0 ac 0.0 PULSE 0 10 20u 0.5u 0.5u 30u 120u 
R_R2 0 2 10k 
R_R3 5 3 1 
V_V2 6 0 dc 10 
R_R1 2 1 10k 
X_U1 3 2 6 4 1 UA741 
V_V3 0 4 dc 10 

*----------------------------------------------

.tran 3e-06 0.0001 0 UIC
.print tran  v(0)
.op

.end
