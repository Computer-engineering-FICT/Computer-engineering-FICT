* /root/laba9/2.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 


*----------------------------------------------

V_V2 7 0 dc 0.0 ac 10meg sin(0.0 10 10000 0 0) 
C_C5 7 5 1e-4 IC=0 
R_R2 2 6 35k 
R_R4 2 3 1k 
.model NPN NPN (is=3.0E-14 NF=1.0 BF=200 IKF=0.5 VAF=100 ISE=7.5E-15 NE=1.4 NR=1.0 BR=4 IKR=0.24 VAR=28 ISC=1.0E-11 NC=1.4 RB=0.1 RE=0.2 RC=0.1 CJC=9.0E-12 MJC=0.35 VJC=0.4 CJE=27.0E-12 TF=0.3E-9 TR=100E-9) 
C_C4 3 4 1e-5 IC=0 
Q_Q1 3 5 1 NPN 
V_V1 2 0 dc 7 
C_C3 4 0 1e-8 IC=0 
C_C2 5 0 1e-7 IC=0 
C_C1 1 0 1e-5 IC=0 
R_R3 1 0 200 
R_R1 6 0 8k 
L_L1 5 4 3.5e-4 

*----------------------------------------------

.ac DEC 10 1 1e+06
.print ac  vm(2)
.op

.end
