* /root/laba1/4.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 

*----------------------------------------------

V_V1 1 0 dc 0.0 ac 0.0 PULSE 0 10 20u 0.5u 0.5u 30u 120u 
C_C1 1 2 0.59n IC=0 
R_R1 2 0 1000 

*----------------------------------------------

.tran 1e-06 0.0001 0 UIC
.print tran  v(1)
.op

.end
