* /root/laba10/1.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/4LB101.model

*----------------------------------------------

.model rmod r (TC1=0 TC2=1e-3) 
R_R3 1 0 10k rmod 
R_R2 3 2 10k  rmod 
R_R1 1 2 10k rmod 
V_V2 0 4 dc 8
V_V1 5 0 dc 8 
X_U1 1 3 5 4 2 4LB101 
C_C1 0 3 4e-3 IC=0 

*----------------------------------------------

.tran 0.0001 0.01 UIC
.print tran  v(1)
.op

.end
