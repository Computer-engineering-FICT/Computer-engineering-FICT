* /root/laba15/4.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/1NPN.model


*----------------------------------------------
.model d d(is=5.72f bv=9.8 rs=7.9 tt=5u cjo=1.67n vj=750m m=504m)
D_D2 3 2 d
R_R1 5 3 2k 
D_D1 3 1 d
V_V1 5 0 dc 0.0 ac 0.0 PULSE 0.0 10 0 0.01u 0.01u 0.5u 1u 
R_R3 2 6 1 
R_R2 4 1 300 
Q_Q1 1 6 0 1NPN 
R_R4 2 0 1k 
V_V2 4 0 dc 10 
vtpi@1 2 6 0 
*----------------------------------------------

.tran 1e-07 5e-06 0 
.print tran  v(4)
.op

.end
