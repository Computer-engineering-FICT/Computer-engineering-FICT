
library IEEE;

use IEEE.STD_LOGIC_1164.all;

entity OR64_SC is
	
	port (D : in STD_LOGIC_VECTOR(63 downto 0); Z : out STD_LOGIC);
	
end OR64_SC;
