

architecture PLM4_DC7 of PLM_4 is
begin
	
	Y <= (D and C and B and A) after td;
	
end PLM4_DC7;