astable
*SPICE_NET
.MODEL QSTD NPN IS=1E-16 BF=50 BR=0.1 RB=50 RC=10 TF=.12NS
+ TR=5NS CJE=0.4PF PE=0.8 ME=0.4 CJC=0.5PF PC=0.8 MC=0.333
+ CCS=1PF VA=50
VIN 6 0 PULSE 0 5 0 1US 1US 100US 100US
Q2 2 5 0 QSTD
Q1 1 3 0 QSTD
C1 1 5 150PF
C2 3 2 150PF
RB1 4 3 30K
RC2 4 2 1K
RC1 4 1 1K
RB2 6 5 30K
VCC 4 0 5
.TRAN 1e-007 10US 0 0
.TEMP 27
.PLOT TRAN V(1) 6,-5
.PLOT TRAN V(2) 6,-5
.PLOT TRAN V(3) 6,-5
.PRINT TRAN V(1) V(2) V(3) 
.END

