* /root/laba7/1.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/UA741.model

*----------------------------------------------

R_R2 3 2 10k 
V_V1 3 0 dc 0 ac 100m sin(0.0 1 10000 0 0) 
R_R1 2 1 10k 
X_U1 0 2 5 4 1 UA741 
V_V2 5 0 dc 10 
V_V3 0 4 dc 10 
VTPI@1 3 2 0
*----------------------------------------------

.dc V_V1 -10 10 1
.print dc   v(3)
.ac DEC 10 1 1e+08
.print ac  vm(3)
.op

.end
