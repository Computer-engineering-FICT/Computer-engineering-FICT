* /root/laba17/1.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 

*----------------------------------------------

V_V2 2 0 dc 5 
R_R1 1 2 500 
V_V1 3 0 dc 0.0 ac 0.0 PULSE 0.0 5 0 0.01u 0.01u 0.2u 1u 
M_M1 1 3 0 0 nmos 
.model nmos nmos (vto=2.5 KP=0.06  gamma=0 phi=600m lambda=35.07m rd=1.10826 rs=187.488m  cgso=300n cgdo=300n cgbo=100n tox=0 nsub=0 tpg=1 uo=600 ) 

*----------------------------------------------

.tran 1e-07 2e-06 0 UIC
.print tran  v(2)
.dc V_V1 0 7 0.1
.print dc   v(2)
.op

.end
