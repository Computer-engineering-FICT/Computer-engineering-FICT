* /root/laba14/2.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/1NPN.model

*----------------------------------------------

V_V3 4 0 dc 0.0 ac 0.0 PULSE 0.0 10 0 0.01u 0.01u 30u 120u 
V_V2 2 0 dc 10 
V_V1 5 0 dc 0.0 ac 0.0 PULSE 0.0 10 0 0.01u 0.01u 30u 120u 
R_R3 1 4 1 
Q_Q1 1 3 0 1NPN 
R_R1 5 3 5k 
R_R2 2 1 400 
vtpi@1 4 1 0
*----------------------------------------------

.dc V_V1 0 10 0.1 V_V3 0 10 0.1
.print dc   v(2)
.op

.end
