UA709
.MODEL QNL NPN BF=80 RB=100 CCS=2PF TF=0.3NS TR=6NS CJE=3PF CJC=2P VA=50
.MODEL QPL PNP BF=10 RB=20 TF=1NS TR=20NS CJE=6PF CJC=4PF VA=50
VIN 3 0 AC 1 SIN 0 0.2 10KHZ 2.5US
VEE 1 0 -15
Q3 30 15 16 QNL
R7 30 15 10K
R8 30 23 10K
RCOMP 23 24 1.5K
R15 20 17 1K
R1 16 12 25K
R2 16 14 25K
Q1 12 2 18 QNL
Q2 14 6 18 QNL
RS2 6 0 1K
RS1 3 2 1K
RF 2 33 100K
Q11 18 4 5 QNL
Q12 8 4 1 QNL
R3 5 1 2.4K
R4 8 7 18K
R5 7 11 3.6K
R9 7 17 10K
Q4 15 14 9 QNL
Q13 13 13 11 QNL
R6 9 13 3K
Q5 15 9 11 QNL
Q6 23 10 11 QNL
Q7 23 12 10 QNL
R14 10 13 3K
CICOMP 12 24 5000PF
Q8 30 23 20 QNL
Q14 22 11 17 QPL
Q15 1 21 33 QPL
Q10 21 22 19 QNL
R12 22 19 10K
R13 19 1 75
COCOMP 33 22 200PF
R10 17 33 30K
R11 30 21 20K
Q9 30 21 33 QNL
VCC 30 0 15
.PROBE
.TRAN 2.5e-006 250US 0 0
.PLOT TRAN V(33) 14.2444,14.2427
.PLOT TRAN V(23) 14.9996,14.9992
.PLOT TRAN V(3) 0.25,-0.25
.PRINT TRAN V(33) V(23) V(3) 
.AC DEC 10 1 1e+010
.TEMP 101
.PLOT AC VM(33) VM(23) VM(3) 1.5,0
.PLOT AC VP(33) VP(23) VP(3) 50,-600
.PRINT AC VM(33)
.PRINT AC VP(33)
.PRINT AC VM(23)
.PRINT AC VP(23)
.PRINT AC VM(3)
.PRINT AC VP(3)
.END


