ttlinv
*SPICE_NET
.MODEL D1 D RS=40 TT=0.1NS CJO=0.9PF
.MODEL QND NPN BF=50 RB=70 RC=40 CCS=2PF TF=0.1NS TR=10NS
+ CJE=0.9PF CJC=1.5PF PC=0.85 VA=50
Q2 3 2 7 QND
Q3 6 3 4 QND
Q5 10 13 5 QND
D1 4 5 D1
D2 10 9 D1
D3 9 0 D1
RB1 11 12 4K
RC3 11 6 100
RC2 11 3 1.4K
RE2 7 0 1K
VCC 11 0 5
VIN 8 0 PULSE 0 3.5 1NS 1NS 1NS 40NS
RS 8 1 50
Q4 5 7 0 QND
RB5 11 13 4K
Q1 2 12 1 QND
.TRAN 1e-009 100NS 0 0
.PLOT TRAN V(3) 6,0
.PLOT TRAN V(5) 4,0
.PRINT TRAN V(3) V(5) 
.dc VIN 0 5 0.05
.TEMP 0
.PLOT DC V(3) 5.5,0.5
.PLOT DC V(5) 4,0
.PRINT DC V(3)
.PRINT DC V(5)
.END

