* /root/laba19/1.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 

.include /usr/X11R6/share/gnome/oregano/models/NPN.model

*----------------------------------------------

.model diode D ( is=5.72393f bv=6.67 rs=4.1 tt=5u cjo=2.02683n vj=750.143m m=504.468m) 
D_D3 0 1 diode 
V_V2 7 0 dc 5 
D_D4 2 8 diode 
V_V3 3 0 dc 5 
R_R5 8 3 1k 
R_R4 7 2 150 
D_D2 0 1 diode 
D_D1 5 1 diode 
R_R2 1 4 1k 
R_R1 5 6 1 
R_R3 4 0 6k 
V_V1 6 0 dc 0.0 ac 0.0 PULSE 0.0 5 0.0 0.01u 0.01u 0.5u 0.7u 
Q_Q1 2 4 0 NPN 
vtpi@1 6 5 0
*----------------------------------------------

.tran 1e-07 6e-06 0 UIC
.print tran  v(4)
.dc V_V1 0 5 0.1
.print dc   v(4)
.op

.end
