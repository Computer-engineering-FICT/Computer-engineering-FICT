
library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity RAM is
	port (
		CLK : in STD_LOGIC; 								-- ���������� 
		WR  : in STD_LOGIC;  							-- ������ ������
		AP  : in STD_LOGIC_VECTOR(13 downto 0);	-- ����� ������ P ��� ������
		AQ  : in STD_LOGIC_VECTOR(13 downto 0);	-- ����� ������ Q ��� ������
		AD  : in STD_LOGIC_VECTOR(13 downto 0);	-- ����� ������ D ��� ������
		P   : out STD_LOGIC_VECTOR(14 downto 0);	-- ������ ������ P
		Q   : in STD_LOGIC_VECTOR (14 downto 0);	-- ������ ������ Q
		D   : out STD_LOGIC_VECTOR(14 downto 0);	-- ������ ������ D
		OE  : in STD_LOGIC								-- ������ ������ ������������ �����
		);
end RAM;

architecture Behavior of RAM is

begin 
	RAMemory: entity work.RAM8 port map
		
end Behavior;