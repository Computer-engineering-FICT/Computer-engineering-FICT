schmitt
*SPICE_NET
.MODEL QSTD NPN IS=1E-16 BF=50 BR=0.1 RB=50 RC=10 TF=0.12NS
+ TR=5NS CJE=0.4PF PE=0.8 ME=0.4 CJC=0.5PF PC=0.8 MC=0.333
+ CCS=1PF VA=50
Q2 2 6 3 QSTD
Q3 0 2 7 QSTD
Q4 0 2 7 QSTD
RIN 4 1 50
R1 5 6 185
RC1 5 0 50
R2 6 8 760
RE 3 8 260
RTH2 7 0 85
RTH1 7 8 125
CLOAD 7 0 5PF
VEE 8 0 -5
V2 4 0 PULSE -1.6 -1.2 10NS 400NS 400NS 100NS 1000NS
RC2 2 0 100
Q1 5 1 3 QSTD
.TRAN 1e-008 1000NS 0 0
.TEMP 27
.PLOT TRAN V(7) -0.8,-2.5
.PLOT TRAN V(5) -0.2,-0.9
.PLOT TRAN V(2) 0,-1.5
.PRINT TRAN V(7) V(5) V(2) 
.END

