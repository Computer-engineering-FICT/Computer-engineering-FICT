
library IEEE;

use IEEE.STD_LOGIC_1164.all;

entity OR8_SC is
	
	port (D : in STD_LOGIC_VECTOR(7 downto 0); Z : out STD_LOGIC);
	
end OR8_SC;
