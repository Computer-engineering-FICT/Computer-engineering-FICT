* /root/laba2/laba2.oregano
*----------------------------------------------
*	NGSPICE - NETLIST
.options NOPAGE 
.include /usr/X11R6/share/gnome/oregano/models/NPN.model

*----------------------------------------------

R_R1 4 2 1k 
V_V1 4 0 dc 0.0 ac 0.0 sin(0.0 5.0 10000 0 0) 
R_R2 1 3 700 
Q_Q1 1 2 0 NPN 
V_V3 3 0 dc 10 
VTPI@1 4 2 0
*----------------------------------------------

.dc V_V1 -1.5 5.5 0.01
.print dc   v(3)
.op

.end
