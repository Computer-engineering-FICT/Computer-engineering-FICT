rca3040
.MODEL QNL NPN BF=80 RB=100 CCS=2PF TF=0.3NS TR=6NS CJE=3PF
+ CJC=2PF VA=50
R6 12 6 1.32K
R7 12 15 4.5K
R8 12 13 1.32K
Q10 12 13 1 QNL
R9 1 0 5.25K
Q11 12 6 2 QNL
R10 2 0 5.25K
VIN 3 0 SIN 0 0.1 50MEG 0.5NS AC 1
RS1 3 4 1K
Q1 12 4 5 QNL
Q3 16 5 8 QNL
R1 5 19 4.8K
Q5 6 15 16 QNL
Q7 15 15 7 QNL
Q8 7 7 0 QNL
Q9 8 10 9 QNL
R3 9 19 811
R4 10 19 2.17K
R5 10 0 820
R2 18 19 4.8K
Q6 13 15 17 QNL
Q4 17 18 8 QNL
VEE 19 0 -15
Q2 12 20 18 QNL
RS2 20 0 1K
VCC 12 0 15
.TRAN 5e-010 50NS 0 0
.PLOT TRAN V(2) V(1) 15,0
.PRINT TRAN V(2) V(1) 
.AC DEC 20 1 1e+010
.PLOT AC VM(2) VM(1) 150,0
.PLOT AC VP(2) VP(1) 250,-600
.PRINT AC VM(2)
.PRINT AC VP(2)
.PRINT AC VM(1)
.PRINT AC VP(1)
.dc VIN -0.25 0.25 0.005
.TEMP 201
.PLOT DC V(2) 20,0
.PRINT DC V(1)
.PRINT DC V(2)
.END

